* Coriolis Structural SPICE Driver
* Generated on Apr 11, 2023, 23:43
* Cell/Subckt "arlet6502_cts_r".
* 
* INTERF we
* INTERF vss
* INTERF vdd
* INTERF reset
* INTERF rdy
* INTERF nmi
* INTERF irq
* INTERF do[7]
* INTERF do[6]
* INTERF do[5]
* INTERF do[4]
* INTERF do[3]
* INTERF do[2]
* INTERF do[1]
* INTERF do[0]
* INTERF di[7]
* INTERF di[6]
* INTERF di[5]
* INTERF di[4]
* INTERF di[3]
* INTERF di[2]
* INTERF di[1]
* INTERF di[0]
* INTERF clk
* INTERF a[9]
* INTERF a[8]
* INTERF a[7]
* INTERF a[6]
* INTERF a[5]
* INTERF a[4]
* INTERF a[3]
* INTERF a[2]
* INTERF a[15]
* INTERF a[14]
* INTERF a[13]
* INTERF a[12]
* INTERF a[11]
* INTERF a[10]
* INTERF a[1]
* INTERF a[0]

* Terminal models (aka standard cells) used througout all the hierarchy.
.include decap_w0.spi
.include o2_x2.spi
.include mx2_x2.spi
.include ao22_x2.spi
.include a3_x2.spi
.include oa22_x2.spi
.include nand3_x0.spi
.include nand2_x0.spi
.include nand4_x0.spi
.include a2_x2.spi
.include sff1_x4.spi
.include tie.spi
.include o4_x2.spi
.include nxr2_x1.spi
.include buf_x4.spi
.include a4_x2.spi
.include nor2_x0.spi
.include mx3_x2.spi
.include inv_x0.spi
.include nor3_x0.spi
.include nor4_x0.spi
.include o3_x2.spi
.include xr2_x1.spi

* Non-terminal models (part of the user's design hierarchy).

.subckt arlet6502_cts_r 0 1 2 8 9 10 177 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 213 1969 1970 1971 1972 1973 1974 1975 1976 1977 1978 1979 1980 1981 1982 1983 1984
* NET     0 = we
* NET     1 = vss
* NET     2 = vdd
* NET     3 = reset_root_tr_0
* NET     4 = reset_root_tl_0
* NET     5 = reset_root_br_0
* NET     6 = reset_root_bl_0
* NET     7 = reset_root_0
* NET     8 = reset
* NET     9 = rdy
* NET    10 = nmi
* NET    11 = mos6502_z
* NET    12 = mos6502_write_back
* NET    13 = mos6502_v
* NET    14 = mos6502_store
* NET    15 = mos6502_state_bit4_hfns_2
* NET    16 = mos6502_state_bit4_hfns_1
* NET    17 = mos6502_state_bit4_hfns_0
* NET    18 = mos6502_state_bit3_hfns_2
* NET    19 = mos6502_state_bit3_hfns_1
* NET    20 = mos6502_state_bit3_hfns_0
* NET    21 = mos6502_state_bit2_hfns_2
* NET    22 = mos6502_state_bit2_hfns_1
* NET    23 = mos6502_state_bit2_hfns_0
* NET    24 = mos6502_state_bit0_hfns_2
* NET    25 = mos6502_state_bit0_hfns_1
* NET    26 = mos6502_state_bit0_hfns_0
* NET    27 = mos6502_state[5]
* NET    28 = mos6502_state[4]
* NET    29 = mos6502_state[3]
* NET    30 = mos6502_state[2]
* NET    31 = mos6502_state[1]
* NET    32 = mos6502_state[0]
* NET    33 = mos6502_src_reg[1]
* NET    34 = mos6502_src_reg[0]
* NET    35 = mos6502_shift_right
* NET    36 = mos6502_shift
* NET    37 = mos6502_sei
* NET    38 = mos6502_sed
* NET    39 = mos6502_sec
* NET    40 = mos6502_rotate
* NET    41 = mos6502_res
* NET    42 = mos6502_plp
* NET    43 = mos6502_php
* NET    44 = mos6502_pc[9]
* NET    45 = mos6502_pc[8]
* NET    46 = mos6502_pc[7]
* NET    47 = mos6502_pc[6]
* NET    48 = mos6502_pc[5]
* NET    49 = mos6502_pc[4]
* NET    50 = mos6502_pc[3]
* NET    51 = mos6502_pc[2]
* NET    52 = mos6502_pc[15]
* NET    53 = mos6502_pc[14]
* NET    54 = mos6502_pc[13]
* NET    55 = mos6502_pc[12]
* NET    56 = mos6502_pc[11]
* NET    57 = mos6502_pc[10]
* NET    58 = mos6502_pc[1]
* NET    59 = mos6502_pc[0]
* NET    60 = mos6502_op[3]
* NET    61 = mos6502_op[2]
* NET    62 = mos6502_op[1]
* NET    63 = mos6502_op[0]
* NET    64 = mos6502_nmi_edge
* NET    65 = mos6502_nmi_1
* NET    66 = mos6502_n
* NET    67 = mos6502_load_reg
* NET    68 = mos6502_load_only
* NET    69 = mos6502_irhold_valid_hfns_2
* NET    70 = mos6502_irhold_valid_hfns_1
* NET    71 = mos6502_irhold_valid_hfns_0
* NET    72 = mos6502_irhold_valid
* NET    73 = mos6502_irhold[7]
* NET    74 = mos6502_irhold[6]
* NET    75 = mos6502_irhold[5]
* NET    76 = mos6502_irhold[4]
* NET    77 = mos6502_irhold[3]
* NET    78 = mos6502_irhold[2]
* NET    79 = mos6502_irhold[1]
* NET    80 = mos6502_irhold[0]
* NET    81 = mos6502_index_y
* NET    82 = mos6502_inc
* NET    83 = mos6502_i
* NET    84 = mos6502_dst_reg[1]
* NET    85 = mos6502_dst_reg[0]
* NET    86 = mos6502_dimux[7]
* NET    87 = mos6502_dimux[6]
* NET    88 = mos6502_dimux[5]
* NET    89 = mos6502_dimux[4]
* NET    90 = mos6502_dimux[3]
* NET    91 = mos6502_dimux[2]
* NET    92 = mos6502_dimux[1]
* NET    93 = mos6502_dimux[0]
* NET    94 = mos6502_dihold[7]
* NET    95 = mos6502_dihold[6]
* NET    96 = mos6502_dihold[5]
* NET    97 = mos6502_dihold[4]
* NET    98 = mos6502_dihold[3]
* NET    99 = mos6502_dihold[2]
* NET   100 = mos6502_dihold[1]
* NET   101 = mos6502_dihold[0]
* NET   102 = mos6502_d
* NET   103 = mos6502_cond_code[2]
* NET   104 = mos6502_cond_code[1]
* NET   105 = mos6502_cond_code[0]
* NET   106 = mos6502_compare
* NET   107 = mos6502_clv
* NET   108 = mos6502_cli
* NET   109 = mos6502_cld
* NET   110 = mos6502_clc
* NET   111 = mos6502_c
* NET   112 = mos6502_bit_ins
* NET   113 = mos6502_backwards
* NET   114 = mos6502_axys_3_7
* NET   115 = mos6502_axys_3_6
* NET   116 = mos6502_axys_3_5
* NET   117 = mos6502_axys_3_4
* NET   118 = mos6502_axys_3_3
* NET   119 = mos6502_axys_3_2
* NET   120 = mos6502_axys_3_1
* NET   121 = mos6502_axys_3_0
* NET   122 = mos6502_axys_2_7
* NET   123 = mos6502_axys_2_6
* NET   124 = mos6502_axys_2_5
* NET   125 = mos6502_axys_2_4
* NET   126 = mos6502_axys_2_3
* NET   127 = mos6502_axys_2_2
* NET   128 = mos6502_axys_2_1
* NET   129 = mos6502_axys_2_0
* NET   130 = mos6502_axys_1_7
* NET   131 = mos6502_axys_1_6
* NET   132 = mos6502_axys_1_5
* NET   133 = mos6502_axys_1_4
* NET   134 = mos6502_axys_1_3
* NET   135 = mos6502_axys_1_2
* NET   136 = mos6502_axys_1_1
* NET   137 = mos6502_axys_1_0
* NET   138 = mos6502_axys_0_7
* NET   139 = mos6502_axys_0_6
* NET   140 = mos6502_axys_0_5
* NET   141 = mos6502_axys_0_4
* NET   142 = mos6502_axys_0_3
* NET   143 = mos6502_axys_0_2
* NET   144 = mos6502_axys_0_1
* NET   145 = mos6502_axys_0_0
* NET   146 = mos6502_alu_out[7]
* NET   147 = mos6502_alu_out[6]
* NET   148 = mos6502_alu_out[5]
* NET   149 = mos6502_alu_out[4]
* NET   150 = mos6502_alu_out[3]
* NET   151 = mos6502_alu_out[2]
* NET   152 = mos6502_alu_out[1]
* NET   153 = mos6502_alu_out[0]
* NET   154 = mos6502_alu_hc
* NET   155 = mos6502_alu_co
* NET   156 = mos6502_alu_bi7
* NET   157 = mos6502_alu_ai7
* NET   158 = mos6502_adj_bcd
* NET   159 = mos6502_adc_sbc
* NET   160 = mos6502_adc_bcd
* NET   161 = mos6502_abl[7]
* NET   162 = mos6502_abl[6]
* NET   163 = mos6502_abl[5]
* NET   164 = mos6502_abl[4]
* NET   165 = mos6502_abl[3]
* NET   166 = mos6502_abl[2]
* NET   167 = mos6502_abl[1]
* NET   168 = mos6502_abl[0]
* NET   169 = mos6502_abh[7]
* NET   170 = mos6502_abh[6]
* NET   171 = mos6502_abh[5]
* NET   172 = mos6502_abh[4]
* NET   173 = mos6502_abh[3]
* NET   174 = mos6502_abh[2]
* NET   175 = mos6502_abh[1]
* NET   176 = mos6502_abh[0]
* NET   177 = irq
* NET   178 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[5]
* NET   179 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[4]
* NET   180 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[3]
* NET   181 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[2]
* NET   182 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[1]
* NET   183 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[0]
* NET   184 = do[7]
* NET   185 = do[6]
* NET   186 = do[5]
* NET   187 = do[4]
* NET   188 = do[3]
* NET   189 = do[2]
* NET   190 = do[1]
* NET   191 = do[0]
* NET   192 = di[7]
* NET   193 = di[6]
* NET   194 = di[5]
* NET   195 = di[4]
* NET   196 = di[3]
* NET   197 = di[2]
* NET   198 = di[1]
* NET   199 = di[0]
* NET   200 = clk_root_tr_2
* NET   201 = clk_root_tr_1
* NET   202 = clk_root_tr_0
* NET   203 = clk_root_tl_2
* NET   204 = clk_root_tl_1
* NET   205 = clk_root_tl_0
* NET   206 = clk_root_br_2
* NET   207 = clk_root_br_1
* NET   208 = clk_root_br_0
* NET   209 = clk_root_bl_2
* NET   210 = clk_root_bl_1
* NET   211 = clk_root_bl_0
* NET   212 = clk_root_0
* NET   213 = clk
* NET   214 = blockagenet
* NET   215 = abc_11873_new_n999
* NET   216 = abc_11873_new_n998
* NET   217 = abc_11873_new_n997
* NET   218 = abc_11873_new_n996
* NET   219 = abc_11873_new_n995
* NET   220 = abc_11873_new_n994
* NET   221 = abc_11873_new_n993
* NET   222 = abc_11873_new_n992
* NET   223 = abc_11873_new_n991
* NET   224 = abc_11873_new_n989
* NET   225 = abc_11873_new_n988
* NET   226 = abc_11873_new_n987
* NET   227 = abc_11873_new_n986
* NET   228 = abc_11873_new_n985
* NET   229 = abc_11873_new_n984
* NET   230 = abc_11873_new_n983
* NET   231 = abc_11873_new_n982
* NET   232 = abc_11873_new_n981
* NET   233 = abc_11873_new_n980
* NET   234 = abc_11873_new_n979
* NET   235 = abc_11873_new_n977
* NET   236 = abc_11873_new_n976
* NET   237 = abc_11873_new_n975
* NET   238 = abc_11873_new_n974
* NET   239 = abc_11873_new_n973
* NET   240 = abc_11873_new_n972
* NET   241 = abc_11873_new_n971
* NET   242 = abc_11873_new_n970
* NET   243 = abc_11873_new_n969
* NET   244 = abc_11873_new_n968
* NET   245 = abc_11873_new_n967
* NET   246 = abc_11873_new_n965
* NET   247 = abc_11873_new_n964
* NET   248 = abc_11873_new_n963
* NET   249 = abc_11873_new_n962
* NET   250 = abc_11873_new_n961
* NET   251 = abc_11873_new_n960
* NET   252 = abc_11873_new_n959
* NET   253 = abc_11873_new_n958
* NET   254 = abc_11873_new_n957
* NET   255 = abc_11873_new_n956
* NET   256 = abc_11873_new_n955
* NET   257 = abc_11873_new_n954
* NET   258 = abc_11873_new_n953
* NET   259 = abc_11873_new_n952
* NET   260 = abc_11873_new_n951
* NET   261 = abc_11873_new_n950
* NET   262 = abc_11873_new_n949
* NET   263 = abc_11873_new_n948
* NET   264 = abc_11873_new_n947
* NET   265 = abc_11873_new_n946
* NET   266 = abc_11873_new_n945
* NET   267 = abc_11873_new_n944
* NET   268 = abc_11873_new_n943
* NET   269 = abc_11873_new_n942
* NET   270 = abc_11873_new_n941
* NET   271 = abc_11873_new_n940
* NET   272 = abc_11873_new_n939
* NET   273 = abc_11873_new_n938
* NET   274 = abc_11873_new_n937
* NET   275 = abc_11873_new_n936
* NET   276 = abc_11873_new_n935
* NET   277 = abc_11873_new_n934
* NET   278 = abc_11873_new_n933
* NET   279 = abc_11873_new_n932
* NET   280 = abc_11873_new_n931
* NET   281 = abc_11873_new_n930
* NET   282 = abc_11873_new_n929
* NET   283 = abc_11873_new_n928
* NET   284 = abc_11873_new_n927
* NET   285 = abc_11873_new_n925
* NET   286 = abc_11873_new_n924
* NET   287 = abc_11873_new_n923
* NET   288 = abc_11873_new_n922
* NET   289 = abc_11873_new_n921
* NET   290 = abc_11873_new_n920
* NET   291 = abc_11873_new_n918
* NET   292 = abc_11873_new_n917
* NET   293 = abc_11873_new_n916
* NET   294 = abc_11873_new_n915
* NET   295 = abc_11873_new_n914
* NET   296 = abc_11873_new_n913
* NET   297 = abc_11873_new_n912
* NET   298 = abc_11873_new_n911
* NET   299 = abc_11873_new_n910
* NET   300 = abc_11873_new_n909
* NET   301 = abc_11873_new_n908
* NET   302 = abc_11873_new_n906
* NET   303 = abc_11873_new_n905
* NET   304 = abc_11873_new_n904
* NET   305 = abc_11873_new_n903
* NET   306 = abc_11873_new_n902
* NET   307 = abc_11873_new_n901
* NET   308 = abc_11873_new_n900
* NET   309 = abc_11873_new_n899
* NET   310 = abc_11873_new_n897
* NET   311 = abc_11873_new_n896
* NET   312 = abc_11873_new_n895
* NET   313 = abc_11873_new_n894
* NET   314 = abc_11873_new_n893
* NET   315 = abc_11873_new_n892
* NET   316 = abc_11873_new_n891
* NET   317 = abc_11873_new_n890
* NET   318 = abc_11873_new_n889
* NET   319 = abc_11873_new_n888
* NET   320 = abc_11873_new_n887
* NET   321 = abc_11873_new_n886
* NET   322 = abc_11873_new_n885
* NET   323 = abc_11873_new_n884
* NET   324 = abc_11873_new_n883
* NET   325 = abc_11873_new_n882
* NET   326 = abc_11873_new_n881
* NET   327 = abc_11873_new_n880
* NET   328 = abc_11873_new_n879
* NET   329 = abc_11873_new_n878
* NET   330 = abc_11873_new_n877
* NET   331 = abc_11873_new_n876
* NET   332 = abc_11873_new_n875
* NET   333 = abc_11873_new_n874
* NET   334 = abc_11873_new_n873
* NET   335 = abc_11873_new_n872
* NET   336 = abc_11873_new_n871
* NET   337 = abc_11873_new_n870
* NET   338 = abc_11873_new_n869
* NET   339 = abc_11873_new_n868
* NET   340 = abc_11873_new_n866
* NET   341 = abc_11873_new_n865
* NET   342 = abc_11873_new_n864
* NET   343 = abc_11873_new_n863
* NET   344 = abc_11873_new_n862
* NET   345 = abc_11873_new_n861
* NET   346 = abc_11873_new_n860
* NET   347 = abc_11873_new_n859
* NET   348 = abc_11873_new_n858
* NET   349 = abc_11873_new_n857
* NET   350 = abc_11873_new_n856
* NET   351 = abc_11873_new_n855
* NET   352 = abc_11873_new_n854
* NET   353 = abc_11873_new_n853
* NET   354 = abc_11873_new_n852
* NET   355 = abc_11873_new_n851
* NET   356 = abc_11873_new_n850
* NET   357 = abc_11873_new_n849
* NET   358 = abc_11873_new_n848
* NET   359 = abc_11873_new_n847
* NET   360 = abc_11873_new_n846
* NET   361 = abc_11873_new_n845
* NET   362 = abc_11873_new_n844
* NET   363 = abc_11873_new_n843
* NET   364 = abc_11873_new_n842
* NET   365 = abc_11873_new_n841
* NET   366 = abc_11873_new_n840
* NET   367 = abc_11873_new_n839
* NET   368 = abc_11873_new_n838
* NET   369 = abc_11873_new_n837
* NET   370 = abc_11873_new_n836
* NET   371 = abc_11873_new_n835
* NET   372 = abc_11873_new_n834
* NET   373 = abc_11873_new_n833
* NET   374 = abc_11873_new_n832
* NET   375 = abc_11873_new_n831
* NET   376 = abc_11873_new_n830
* NET   377 = abc_11873_new_n829
* NET   378 = abc_11873_new_n828
* NET   379 = abc_11873_new_n827
* NET   380 = abc_11873_new_n826
* NET   381 = abc_11873_new_n825
* NET   382 = abc_11873_new_n824
* NET   383 = abc_11873_new_n823
* NET   384 = abc_11873_new_n822
* NET   385 = abc_11873_new_n821
* NET   386 = abc_11873_new_n820
* NET   387 = abc_11873_new_n819
* NET   388 = abc_11873_new_n818
* NET   389 = abc_11873_new_n817
* NET   390 = abc_11873_new_n816
* NET   391 = abc_11873_new_n814
* NET   392 = abc_11873_new_n813
* NET   393 = abc_11873_new_n812
* NET   394 = abc_11873_new_n811
* NET   395 = abc_11873_new_n810
* NET   396 = abc_11873_new_n809
* NET   397 = abc_11873_new_n808
* NET   398 = abc_11873_new_n807
* NET   399 = abc_11873_new_n806
* NET   400 = abc_11873_new_n805
* NET   401 = abc_11873_new_n804
* NET   402 = abc_11873_new_n803
* NET   403 = abc_11873_new_n802
* NET   404 = abc_11873_new_n801
* NET   405 = abc_11873_new_n800
* NET   406 = abc_11873_new_n799
* NET   407 = abc_11873_new_n798
* NET   408 = abc_11873_new_n797
* NET   409 = abc_11873_new_n796
* NET   410 = abc_11873_new_n795
* NET   411 = abc_11873_new_n794
* NET   412 = abc_11873_new_n793
* NET   413 = abc_11873_new_n792
* NET   414 = abc_11873_new_n791
* NET   415 = abc_11873_new_n790
* NET   416 = abc_11873_new_n789
* NET   417 = abc_11873_new_n788
* NET   418 = abc_11873_new_n787
* NET   419 = abc_11873_new_n786
* NET   420 = abc_11873_new_n785
* NET   421 = abc_11873_new_n784
* NET   422 = abc_11873_new_n783
* NET   423 = abc_11873_new_n782
* NET   424 = abc_11873_new_n781
* NET   425 = abc_11873_new_n780
* NET   426 = abc_11873_new_n779
* NET   427 = abc_11873_new_n778
* NET   428 = abc_11873_new_n777
* NET   429 = abc_11873_new_n776
* NET   430 = abc_11873_new_n775
* NET   431 = abc_11873_new_n774
* NET   432 = abc_11873_new_n773
* NET   433 = abc_11873_new_n772
* NET   434 = abc_11873_new_n771
* NET   435 = abc_11873_new_n770
* NET   436 = abc_11873_new_n769
* NET   437 = abc_11873_new_n768
* NET   438 = abc_11873_new_n767
* NET   439 = abc_11873_new_n766
* NET   440 = abc_11873_new_n765
* NET   441 = abc_11873_new_n764
* NET   442 = abc_11873_new_n763
* NET   443 = abc_11873_new_n762
* NET   444 = abc_11873_new_n761
* NET   445 = abc_11873_new_n760
* NET   446 = abc_11873_new_n759
* NET   447 = abc_11873_new_n758
* NET   448 = abc_11873_new_n757
* NET   449 = abc_11873_new_n756
* NET   450 = abc_11873_new_n755
* NET   451 = abc_11873_new_n754
* NET   452 = abc_11873_new_n753
* NET   453 = abc_11873_new_n752
* NET   454 = abc_11873_new_n751
* NET   455 = abc_11873_new_n750
* NET   456 = abc_11873_new_n749
* NET   457 = abc_11873_new_n748
* NET   458 = abc_11873_new_n747
* NET   459 = abc_11873_new_n746
* NET   460 = abc_11873_new_n745
* NET   461 = abc_11873_new_n744
* NET   462 = abc_11873_new_n743
* NET   463 = abc_11873_new_n742
* NET   464 = abc_11873_new_n740
* NET   465 = abc_11873_new_n739
* NET   466 = abc_11873_new_n738
* NET   467 = abc_11873_new_n737
* NET   468 = abc_11873_new_n736
* NET   469 = abc_11873_new_n735
* NET   470 = abc_11873_new_n734
* NET   471 = abc_11873_new_n733
* NET   472 = abc_11873_new_n732
* NET   473 = abc_11873_new_n731
* NET   474 = abc_11873_new_n730
* NET   475 = abc_11873_new_n729
* NET   476 = abc_11873_new_n728
* NET   477 = abc_11873_new_n727
* NET   478 = abc_11873_new_n726
* NET   479 = abc_11873_new_n725
* NET   480 = abc_11873_new_n724
* NET   481 = abc_11873_new_n723
* NET   482 = abc_11873_new_n722
* NET   483 = abc_11873_new_n721
* NET   484 = abc_11873_new_n720
* NET   485 = abc_11873_new_n719
* NET   486 = abc_11873_new_n718
* NET   487 = abc_11873_new_n717
* NET   488 = abc_11873_new_n716
* NET   489 = abc_11873_new_n715
* NET   490 = abc_11873_new_n714
* NET   491 = abc_11873_new_n713
* NET   492 = abc_11873_new_n712
* NET   493 = abc_11873_new_n711
* NET   494 = abc_11873_new_n710
* NET   495 = abc_11873_new_n709
* NET   496 = abc_11873_new_n708
* NET   497 = abc_11873_new_n707
* NET   498 = abc_11873_new_n706
* NET   499 = abc_11873_new_n705
* NET   500 = abc_11873_new_n704
* NET   501 = abc_11873_new_n703
* NET   502 = abc_11873_new_n702
* NET   503 = abc_11873_new_n701
* NET   504 = abc_11873_new_n700
* NET   505 = abc_11873_new_n699
* NET   506 = abc_11873_new_n698
* NET   507 = abc_11873_new_n697
* NET   508 = abc_11873_new_n696
* NET   509 = abc_11873_new_n695
* NET   510 = abc_11873_new_n694
* NET   511 = abc_11873_new_n693
* NET   512 = abc_11873_new_n692
* NET   513 = abc_11873_new_n691
* NET   514 = abc_11873_new_n690
* NET   515 = abc_11873_new_n689
* NET   516 = abc_11873_new_n688
* NET   517 = abc_11873_new_n687
* NET   518 = abc_11873_new_n686
* NET   519 = abc_11873_new_n685
* NET   520 = abc_11873_new_n684
* NET   521 = abc_11873_new_n683
* NET   522 = abc_11873_new_n682
* NET   523 = abc_11873_new_n681
* NET   524 = abc_11873_new_n680
* NET   525 = abc_11873_new_n679
* NET   526 = abc_11873_new_n678
* NET   527 = abc_11873_new_n677
* NET   528 = abc_11873_new_n676
* NET   529 = abc_11873_new_n675
* NET   530 = abc_11873_new_n674
* NET   531 = abc_11873_new_n673
* NET   532 = abc_11873_new_n672
* NET   533 = abc_11873_new_n671
* NET   534 = abc_11873_new_n670
* NET   535 = abc_11873_new_n669
* NET   536 = abc_11873_new_n668
* NET   537 = abc_11873_new_n667
* NET   538 = abc_11873_new_n666
* NET   539 = abc_11873_new_n665
* NET   540 = abc_11873_new_n664
* NET   541 = abc_11873_new_n663
* NET   542 = abc_11873_new_n662
* NET   543 = abc_11873_new_n661
* NET   544 = abc_11873_new_n660
* NET   545 = abc_11873_new_n659
* NET   546 = abc_11873_new_n658
* NET   547 = abc_11873_new_n657
* NET   548 = abc_11873_new_n656_hfns_2
* NET   549 = abc_11873_new_n656_hfns_1
* NET   550 = abc_11873_new_n656_hfns_0
* NET   551 = abc_11873_new_n656
* NET   552 = abc_11873_new_n655
* NET   553 = abc_11873_new_n654
* NET   554 = abc_11873_new_n653
* NET   555 = abc_11873_new_n652
* NET   556 = abc_11873_new_n651
* NET   557 = abc_11873_new_n650
* NET   558 = abc_11873_new_n649
* NET   559 = abc_11873_new_n648
* NET   560 = abc_11873_new_n647
* NET   561 = abc_11873_new_n646
* NET   562 = abc_11873_new_n645
* NET   563 = abc_11873_new_n644
* NET   564 = abc_11873_new_n643
* NET   565 = abc_11873_new_n642
* NET   566 = abc_11873_new_n641
* NET   567 = abc_11873_new_n640
* NET   568 = abc_11873_new_n639
* NET   569 = abc_11873_new_n638
* NET   570 = abc_11873_new_n637
* NET   571 = abc_11873_new_n636
* NET   572 = abc_11873_new_n635
* NET   573 = abc_11873_new_n634
* NET   574 = abc_11873_new_n633
* NET   575 = abc_11873_new_n632
* NET   576 = abc_11873_new_n631
* NET   577 = abc_11873_new_n630
* NET   578 = abc_11873_new_n629
* NET   579 = abc_11873_new_n628
* NET   580 = abc_11873_new_n627
* NET   581 = abc_11873_new_n626
* NET   582 = abc_11873_new_n625
* NET   583 = abc_11873_new_n624
* NET   584 = abc_11873_new_n623
* NET   585 = abc_11873_new_n622
* NET   586 = abc_11873_new_n621
* NET   587 = abc_11873_new_n620
* NET   588 = abc_11873_new_n619
* NET   589 = abc_11873_new_n618
* NET   590 = abc_11873_new_n617
* NET   591 = abc_11873_new_n616
* NET   592 = abc_11873_new_n615
* NET   593 = abc_11873_new_n614
* NET   594 = abc_11873_new_n613
* NET   595 = abc_11873_new_n612
* NET   596 = abc_11873_new_n611
* NET   597 = abc_11873_new_n610
* NET   598 = abc_11873_new_n609
* NET   599 = abc_11873_new_n608
* NET   600 = abc_11873_new_n607
* NET   601 = abc_11873_new_n606
* NET   602 = abc_11873_new_n605
* NET   603 = abc_11873_new_n604
* NET   604 = abc_11873_new_n603
* NET   605 = abc_11873_new_n602
* NET   606 = abc_11873_new_n601
* NET   607 = abc_11873_new_n600
* NET   608 = abc_11873_new_n599
* NET   609 = abc_11873_new_n598
* NET   610 = abc_11873_new_n597
* NET   611 = abc_11873_new_n596
* NET   612 = abc_11873_new_n595
* NET   613 = abc_11873_new_n594
* NET   614 = abc_11873_new_n593
* NET   615 = abc_11873_new_n592
* NET   616 = abc_11873_new_n591
* NET   617 = abc_11873_new_n590
* NET   618 = abc_11873_new_n589
* NET   619 = abc_11873_new_n588
* NET   620 = abc_11873_new_n587
* NET   621 = abc_11873_new_n586
* NET   622 = abc_11873_new_n585
* NET   623 = abc_11873_new_n584
* NET   624 = abc_11873_new_n583
* NET   625 = abc_11873_new_n582
* NET   626 = abc_11873_new_n581
* NET   627 = abc_11873_new_n580
* NET   628 = abc_11873_new_n579
* NET   629 = abc_11873_new_n578
* NET   630 = abc_11873_new_n577
* NET   631 = abc_11873_new_n576
* NET   632 = abc_11873_new_n575
* NET   633 = abc_11873_new_n574
* NET   634 = abc_11873_new_n573
* NET   635 = abc_11873_new_n572
* NET   636 = abc_11873_new_n571
* NET   637 = abc_11873_new_n570
* NET   638 = abc_11873_new_n569
* NET   639 = abc_11873_new_n568
* NET   640 = abc_11873_new_n567
* NET   641 = abc_11873_new_n566
* NET   642 = abc_11873_new_n565
* NET   643 = abc_11873_new_n564
* NET   644 = abc_11873_new_n563
* NET   645 = abc_11873_new_n562
* NET   646 = abc_11873_new_n561_hfns_2
* NET   647 = abc_11873_new_n561_hfns_1
* NET   648 = abc_11873_new_n561_hfns_0
* NET   649 = abc_11873_new_n561
* NET   650 = abc_11873_new_n560
* NET   651 = abc_11873_new_n559
* NET   652 = abc_11873_new_n558
* NET   653 = abc_11873_new_n557
* NET   654 = abc_11873_new_n556
* NET   655 = abc_11873_new_n555
* NET   656 = abc_11873_new_n554
* NET   657 = abc_11873_new_n553
* NET   658 = abc_11873_new_n552
* NET   659 = abc_11873_new_n551
* NET   660 = abc_11873_new_n550
* NET   661 = abc_11873_new_n549
* NET   662 = abc_11873_new_n548
* NET   663 = abc_11873_new_n547
* NET   664 = abc_11873_new_n546
* NET   665 = abc_11873_new_n545
* NET   666 = abc_11873_new_n544
* NET   667 = abc_11873_new_n543
* NET   668 = abc_11873_new_n542
* NET   669 = abc_11873_new_n541
* NET   670 = abc_11873_new_n540
* NET   671 = abc_11873_new_n539
* NET   672 = abc_11873_new_n538
* NET   673 = abc_11873_new_n537
* NET   674 = abc_11873_new_n536
* NET   675 = abc_11873_new_n535
* NET   676 = abc_11873_new_n534
* NET   677 = abc_11873_new_n533
* NET   678 = abc_11873_new_n532_hfns_3
* NET   679 = abc_11873_new_n532_hfns_2
* NET   680 = abc_11873_new_n532_hfns_1
* NET   681 = abc_11873_new_n532_hfns_0
* NET   682 = abc_11873_new_n532
* NET   683 = abc_11873_new_n531
* NET   684 = abc_11873_new_n530
* NET   685 = abc_11873_new_n529
* NET   686 = abc_11873_new_n528
* NET   687 = abc_11873_new_n527
* NET   688 = abc_11873_new_n526
* NET   689 = abc_11873_new_n525
* NET   690 = abc_11873_new_n524
* NET   691 = abc_11873_new_n523
* NET   692 = abc_11873_new_n522
* NET   693 = abc_11873_new_n521
* NET   694 = abc_11873_new_n520
* NET   695 = abc_11873_new_n519
* NET   696 = abc_11873_new_n518_hfns_2
* NET   697 = abc_11873_new_n518_hfns_1
* NET   698 = abc_11873_new_n518_hfns_0
* NET   699 = abc_11873_new_n518
* NET   700 = abc_11873_new_n517
* NET   701 = abc_11873_new_n516
* NET   702 = abc_11873_new_n515
* NET   703 = abc_11873_new_n514
* NET   704 = abc_11873_new_n513
* NET   705 = abc_11873_new_n512
* NET   706 = abc_11873_new_n511
* NET   707 = abc_11873_new_n510
* NET   708 = abc_11873_new_n509
* NET   709 = abc_11873_new_n508
* NET   710 = abc_11873_new_n507
* NET   711 = abc_11873_new_n506_hfns_2
* NET   712 = abc_11873_new_n506_hfns_1
* NET   713 = abc_11873_new_n506_hfns_0
* NET   714 = abc_11873_new_n506
* NET   715 = abc_11873_new_n505
* NET   716 = abc_11873_new_n504_hfns_3
* NET   717 = abc_11873_new_n504_hfns_2
* NET   718 = abc_11873_new_n504_hfns_1
* NET   719 = abc_11873_new_n504_hfns_0
* NET   720 = abc_11873_new_n504
* NET   721 = abc_11873_new_n503
* NET   722 = abc_11873_new_n502
* NET   723 = abc_11873_new_n501
* NET   724 = abc_11873_new_n500
* NET   725 = abc_11873_new_n499
* NET   726 = abc_11873_new_n498
* NET   727 = abc_11873_new_n497
* NET   728 = abc_11873_new_n496
* NET   729 = abc_11873_new_n495
* NET   730 = abc_11873_new_n494
* NET   731 = abc_11873_new_n493
* NET   732 = abc_11873_new_n492
* NET   733 = abc_11873_new_n491
* NET   734 = abc_11873_new_n490
* NET   735 = abc_11873_new_n489
* NET   736 = abc_11873_new_n488
* NET   737 = abc_11873_new_n487
* NET   738 = abc_11873_new_n486
* NET   739 = abc_11873_new_n485
* NET   740 = abc_11873_new_n484
* NET   741 = abc_11873_new_n483
* NET   742 = abc_11873_new_n482
* NET   743 = abc_11873_new_n481
* NET   744 = abc_11873_new_n480
* NET   745 = abc_11873_new_n479_hfns_2
* NET   746 = abc_11873_new_n479_hfns_1
* NET   747 = abc_11873_new_n479_hfns_0
* NET   748 = abc_11873_new_n479
* NET   749 = abc_11873_new_n478
* NET   750 = abc_11873_new_n477
* NET   751 = abc_11873_new_n476
* NET   752 = abc_11873_new_n475
* NET   753 = abc_11873_new_n474
* NET   754 = abc_11873_new_n473
* NET   755 = abc_11873_new_n472
* NET   756 = abc_11873_new_n471
* NET   757 = abc_11873_new_n470
* NET   758 = abc_11873_new_n469
* NET   759 = abc_11873_new_n468
* NET   760 = abc_11873_new_n467
* NET   761 = abc_11873_new_n466
* NET   762 = abc_11873_new_n465
* NET   763 = abc_11873_new_n464
* NET   764 = abc_11873_new_n463
* NET   765 = abc_11873_new_n462
* NET   766 = abc_11873_new_n461
* NET   767 = abc_11873_new_n460
* NET   768 = abc_11873_new_n459
* NET   769 = abc_11873_new_n458
* NET   770 = abc_11873_new_n457
* NET   771 = abc_11873_new_n456
* NET   772 = abc_11873_new_n455
* NET   773 = abc_11873_new_n454
* NET   774 = abc_11873_new_n453
* NET   775 = abc_11873_new_n452
* NET   776 = abc_11873_new_n451
* NET   777 = abc_11873_new_n450
* NET   778 = abc_11873_new_n449_hfns_2
* NET   779 = abc_11873_new_n449_hfns_1
* NET   780 = abc_11873_new_n449_hfns_0
* NET   781 = abc_11873_new_n449
* NET   782 = abc_11873_new_n448_hfns_2
* NET   783 = abc_11873_new_n448_hfns_1
* NET   784 = abc_11873_new_n448_hfns_0
* NET   785 = abc_11873_new_n448
* NET   786 = abc_11873_new_n447_hfns_2
* NET   787 = abc_11873_new_n447_hfns_1
* NET   788 = abc_11873_new_n447_hfns_0
* NET   789 = abc_11873_new_n447
* NET   790 = abc_11873_new_n446
* NET   791 = abc_11873_new_n445_hfns_4
* NET   792 = abc_11873_new_n445_hfns_3
* NET   793 = abc_11873_new_n445_hfns_2
* NET   794 = abc_11873_new_n445_hfns_1
* NET   795 = abc_11873_new_n445_hfns_0
* NET   796 = abc_11873_new_n445
* NET   797 = abc_11873_new_n444
* NET   798 = abc_11873_new_n443_hfns_2
* NET   799 = abc_11873_new_n443_hfns_1
* NET   800 = abc_11873_new_n443_hfns_0
* NET   801 = abc_11873_new_n443
* NET   802 = abc_11873_new_n441
* NET   803 = abc_11873_new_n439
* NET   804 = abc_11873_new_n437
* NET   805 = abc_11873_new_n435
* NET   806 = abc_11873_new_n433
* NET   807 = abc_11873_new_n431
* NET   808 = abc_11873_new_n429
* NET   809 = abc_11873_new_n427
* NET   810 = abc_11873_new_n426
* NET   811 = abc_11873_new_n425
* NET   812 = abc_11873_new_n424
* NET   813 = abc_11873_new_n423
* NET   814 = abc_11873_new_n422
* NET   815 = abc_11873_new_n421
* NET   816 = abc_11873_new_n420
* NET   817 = abc_11873_new_n419
* NET   818 = abc_11873_new_n418
* NET   819 = abc_11873_new_n417
* NET   820 = abc_11873_new_n416
* NET   821 = abc_11873_new_n415
* NET   822 = abc_11873_new_n414
* NET   823 = abc_11873_new_n413
* NET   824 = abc_11873_new_n412
* NET   825 = abc_11873_new_n411
* NET   826 = abc_11873_new_n410
* NET   827 = abc_11873_new_n409
* NET   828 = abc_11873_new_n408
* NET   829 = abc_11873_new_n407
* NET   830 = abc_11873_new_n406
* NET   831 = abc_11873_new_n405
* NET   832 = abc_11873_new_n404
* NET   833 = abc_11873_new_n403
* NET   834 = abc_11873_new_n402
* NET   835 = abc_11873_new_n401
* NET   836 = abc_11873_new_n400
* NET   837 = abc_11873_new_n399
* NET   838 = abc_11873_new_n398
* NET   839 = abc_11873_new_n397
* NET   840 = abc_11873_new_n396
* NET   841 = abc_11873_new_n395
* NET   842 = abc_11873_new_n394
* NET   843 = abc_11873_new_n393
* NET   844 = abc_11873_new_n392
* NET   845 = abc_11873_new_n391
* NET   846 = abc_11873_new_n390
* NET   847 = abc_11873_new_n389
* NET   848 = abc_11873_new_n388
* NET   849 = abc_11873_new_n387
* NET   850 = abc_11873_new_n386
* NET   851 = abc_11873_new_n385
* NET   852 = abc_11873_new_n384
* NET   853 = abc_11873_new_n383
* NET   854 = abc_11873_new_n382
* NET   855 = abc_11873_new_n381
* NET   856 = abc_11873_new_n380
* NET   857 = abc_11873_new_n379
* NET   858 = abc_11873_new_n378
* NET   859 = abc_11873_new_n377
* NET   860 = abc_11873_new_n376
* NET   861 = abc_11873_new_n375
* NET   862 = abc_11873_new_n374
* NET   863 = abc_11873_new_n373
* NET   864 = abc_11873_new_n372
* NET   865 = abc_11873_new_n371
* NET   866 = abc_11873_new_n370
* NET   867 = abc_11873_new_n369
* NET   868 = abc_11873_new_n368
* NET   869 = abc_11873_new_n367
* NET   870 = abc_11873_new_n366
* NET   871 = abc_11873_new_n365
* NET   872 = abc_11873_new_n364
* NET   873 = abc_11873_new_n363
* NET   874 = abc_11873_new_n362
* NET   875 = abc_11873_new_n361
* NET   876 = abc_11873_new_n360
* NET   877 = abc_11873_new_n359
* NET   878 = abc_11873_new_n358
* NET   879 = abc_11873_new_n357
* NET   880 = abc_11873_new_n356
* NET   881 = abc_11873_new_n355
* NET   882 = abc_11873_new_n354
* NET   883 = abc_11873_new_n353
* NET   884 = abc_11873_new_n352
* NET   885 = abc_11873_new_n351
* NET   886 = abc_11873_new_n350
* NET   887 = abc_11873_new_n349
* NET   888 = abc_11873_new_n348
* NET   889 = abc_11873_new_n347
* NET   890 = abc_11873_new_n346
* NET   891 = abc_11873_new_n345
* NET   892 = abc_11873_new_n344
* NET   893 = abc_11873_new_n343
* NET   894 = abc_11873_new_n342
* NET   895 = abc_11873_new_n341
* NET   896 = abc_11873_new_n340
* NET   897 = abc_11873_new_n339
* NET   898 = abc_11873_new_n338
* NET   899 = abc_11873_new_n337
* NET   900 = abc_11873_new_n336
* NET   901 = abc_11873_new_n335_hfns_3
* NET   902 = abc_11873_new_n335_hfns_2
* NET   903 = abc_11873_new_n335_hfns_1
* NET   904 = abc_11873_new_n335_hfns_0
* NET   905 = abc_11873_new_n335
* NET   906 = abc_11873_new_n334
* NET   907 = abc_11873_new_n333
* NET   908 = abc_11873_new_n332
* NET   909 = abc_11873_new_n331
* NET   910 = abc_11873_new_n330
* NET   911 = abc_11873_new_n329
* NET   912 = abc_11873_new_n328
* NET   913 = abc_11873_new_n327
* NET   914 = abc_11873_new_n326
* NET   915 = abc_11873_new_n325
* NET   916 = abc_11873_new_n324
* NET   917 = abc_11873_new_n323
* NET   918 = abc_11873_new_n2069
* NET   919 = abc_11873_new_n2068
* NET   920 = abc_11873_new_n2063
* NET   921 = abc_11873_new_n2058
* NET   922 = abc_11873_new_n2057
* NET   923 = abc_11873_new_n2055
* NET   924 = abc_11873_new_n2054
* NET   925 = abc_11873_new_n2053
* NET   926 = abc_11873_new_n2052
* NET   927 = abc_11873_new_n2051
* NET   928 = abc_11873_new_n2050
* NET   929 = abc_11873_new_n2049
* NET   930 = abc_11873_new_n2048
* NET   931 = abc_11873_new_n2047
* NET   932 = abc_11873_new_n2046
* NET   933 = abc_11873_new_n2045
* NET   934 = abc_11873_new_n2044
* NET   935 = abc_11873_new_n2043
* NET   936 = abc_11873_new_n2042
* NET   937 = abc_11873_new_n2041
* NET   938 = abc_11873_new_n2040
* NET   939 = abc_11873_new_n2039
* NET   940 = abc_11873_new_n2038
* NET   941 = abc_11873_new_n2037
* NET   942 = abc_11873_new_n2036
* NET   943 = abc_11873_new_n2035
* NET   944 = abc_11873_new_n2034
* NET   945 = abc_11873_new_n2033
* NET   946 = abc_11873_new_n2032
* NET   947 = abc_11873_new_n2031
* NET   948 = abc_11873_new_n2030
* NET   949 = abc_11873_new_n2029
* NET   950 = abc_11873_new_n2028
* NET   951 = abc_11873_new_n2027
* NET   952 = abc_11873_new_n2026
* NET   953 = abc_11873_new_n2025
* NET   954 = abc_11873_new_n2024
* NET   955 = abc_11873_new_n2023
* NET   956 = abc_11873_new_n2022
* NET   957 = abc_11873_new_n2021
* NET   958 = abc_11873_new_n2020
* NET   959 = abc_11873_new_n2019
* NET   960 = abc_11873_new_n2018
* NET   961 = abc_11873_new_n2017
* NET   962 = abc_11873_new_n2016
* NET   963 = abc_11873_new_n2015
* NET   964 = abc_11873_new_n2014
* NET   965 = abc_11873_new_n2013
* NET   966 = abc_11873_new_n2012
* NET   967 = abc_11873_new_n2011
* NET   968 = abc_11873_new_n2010
* NET   969 = abc_11873_new_n2009
* NET   970 = abc_11873_new_n2008
* NET   971 = abc_11873_new_n2007
* NET   972 = abc_11873_new_n2006
* NET   973 = abc_11873_new_n2005
* NET   974 = abc_11873_new_n2004
* NET   975 = abc_11873_new_n2003
* NET   976 = abc_11873_new_n2002
* NET   977 = abc_11873_new_n2001
* NET   978 = abc_11873_new_n2000
* NET   979 = abc_11873_new_n1999
* NET   980 = abc_11873_new_n1998
* NET   981 = abc_11873_new_n1997
* NET   982 = abc_11873_new_n1996
* NET   983 = abc_11873_new_n1995
* NET   984 = abc_11873_new_n1994
* NET   985 = abc_11873_new_n1993
* NET   986 = abc_11873_new_n1992
* NET   987 = abc_11873_new_n1991
* NET   988 = abc_11873_new_n1990
* NET   989 = abc_11873_new_n1989
* NET   990 = abc_11873_new_n1988
* NET   991 = abc_11873_new_n1987
* NET   992 = abc_11873_new_n1986
* NET   993 = abc_11873_new_n1985
* NET   994 = abc_11873_new_n1984
* NET   995 = abc_11873_new_n1983
* NET   996 = abc_11873_new_n1982
* NET   997 = abc_11873_new_n1981
* NET   998 = abc_11873_new_n1980
* NET   999 = abc_11873_new_n1979
* NET  1000 = abc_11873_new_n1978
* NET  1001 = abc_11873_new_n1977
* NET  1002 = abc_11873_new_n1976
* NET  1003 = abc_11873_new_n1975
* NET  1004 = abc_11873_new_n1974
* NET  1005 = abc_11873_new_n1973
* NET  1006 = abc_11873_new_n1972
* NET  1007 = abc_11873_new_n1971
* NET  1008 = abc_11873_new_n1970
* NET  1009 = abc_11873_new_n1969
* NET  1010 = abc_11873_new_n1968
* NET  1011 = abc_11873_new_n1967
* NET  1012 = abc_11873_new_n1966
* NET  1013 = abc_11873_new_n1965
* NET  1014 = abc_11873_new_n1964
* NET  1015 = abc_11873_new_n1963
* NET  1016 = abc_11873_new_n1962
* NET  1017 = abc_11873_new_n1961
* NET  1018 = abc_11873_new_n1960
* NET  1019 = abc_11873_new_n1959
* NET  1020 = abc_11873_new_n1958
* NET  1021 = abc_11873_new_n1957
* NET  1022 = abc_11873_new_n1956
* NET  1023 = abc_11873_new_n1955
* NET  1024 = abc_11873_new_n1954
* NET  1025 = abc_11873_new_n1953
* NET  1026 = abc_11873_new_n1952
* NET  1027 = abc_11873_new_n1951
* NET  1028 = abc_11873_new_n1950
* NET  1029 = abc_11873_new_n1949
* NET  1030 = abc_11873_new_n1948
* NET  1031 = abc_11873_new_n1947
* NET  1032 = abc_11873_new_n1946
* NET  1033 = abc_11873_new_n1945
* NET  1034 = abc_11873_new_n1944
* NET  1035 = abc_11873_new_n1943
* NET  1036 = abc_11873_new_n1942
* NET  1037 = abc_11873_new_n1941
* NET  1038 = abc_11873_new_n1940
* NET  1039 = abc_11873_new_n1939
* NET  1040 = abc_11873_new_n1938
* NET  1041 = abc_11873_new_n1937
* NET  1042 = abc_11873_new_n1936
* NET  1043 = abc_11873_new_n1935
* NET  1044 = abc_11873_new_n1934
* NET  1045 = abc_11873_new_n1933
* NET  1046 = abc_11873_new_n1932
* NET  1047 = abc_11873_new_n1931
* NET  1048 = abc_11873_new_n1930
* NET  1049 = abc_11873_new_n1929
* NET  1050 = abc_11873_new_n1928
* NET  1051 = abc_11873_new_n1927
* NET  1052 = abc_11873_new_n1926
* NET  1053 = abc_11873_new_n1925
* NET  1054 = abc_11873_new_n1924
* NET  1055 = abc_11873_new_n1923
* NET  1056 = abc_11873_new_n1922
* NET  1057 = abc_11873_new_n1921
* NET  1058 = abc_11873_new_n1920
* NET  1059 = abc_11873_new_n1919
* NET  1060 = abc_11873_new_n1918
* NET  1061 = abc_11873_new_n1917
* NET  1062 = abc_11873_new_n1916
* NET  1063 = abc_11873_new_n1915
* NET  1064 = abc_11873_new_n1914
* NET  1065 = abc_11873_new_n1913
* NET  1066 = abc_11873_new_n1912
* NET  1067 = abc_11873_new_n1911
* NET  1068 = abc_11873_new_n1910
* NET  1069 = abc_11873_new_n1909
* NET  1070 = abc_11873_new_n1908
* NET  1071 = abc_11873_new_n1907
* NET  1072 = abc_11873_new_n1906
* NET  1073 = abc_11873_new_n1905
* NET  1074 = abc_11873_new_n1904
* NET  1075 = abc_11873_new_n1903
* NET  1076 = abc_11873_new_n1902
* NET  1077 = abc_11873_new_n1901
* NET  1078 = abc_11873_new_n1900
* NET  1079 = abc_11873_new_n1899
* NET  1080 = abc_11873_new_n1898
* NET  1081 = abc_11873_new_n1897
* NET  1082 = abc_11873_new_n1896
* NET  1083 = abc_11873_new_n1895
* NET  1084 = abc_11873_new_n1894
* NET  1085 = abc_11873_new_n1893
* NET  1086 = abc_11873_new_n1892
* NET  1087 = abc_11873_new_n1891
* NET  1088 = abc_11873_new_n1890
* NET  1089 = abc_11873_new_n1889
* NET  1090 = abc_11873_new_n1888
* NET  1091 = abc_11873_new_n1887
* NET  1092 = abc_11873_new_n1886
* NET  1093 = abc_11873_new_n1885
* NET  1094 = abc_11873_new_n1884
* NET  1095 = abc_11873_new_n1883
* NET  1096 = abc_11873_new_n1882
* NET  1097 = abc_11873_new_n1881
* NET  1098 = abc_11873_new_n1880
* NET  1099 = abc_11873_new_n1879
* NET  1100 = abc_11873_new_n1878
* NET  1101 = abc_11873_new_n1877
* NET  1102 = abc_11873_new_n1876
* NET  1103 = abc_11873_new_n1875
* NET  1104 = abc_11873_new_n1874
* NET  1105 = abc_11873_new_n1873
* NET  1106 = abc_11873_new_n1872
* NET  1107 = abc_11873_new_n1871
* NET  1108 = abc_11873_new_n1870
* NET  1109 = abc_11873_new_n1869
* NET  1110 = abc_11873_new_n1868
* NET  1111 = abc_11873_new_n1867
* NET  1112 = abc_11873_new_n1866
* NET  1113 = abc_11873_new_n1865
* NET  1114 = abc_11873_new_n1864
* NET  1115 = abc_11873_new_n1863
* NET  1116 = abc_11873_new_n1862
* NET  1117 = abc_11873_new_n1861
* NET  1118 = abc_11873_new_n1860
* NET  1119 = abc_11873_new_n1859
* NET  1120 = abc_11873_new_n1858
* NET  1121 = abc_11873_new_n1857
* NET  1122 = abc_11873_new_n1856
* NET  1123 = abc_11873_new_n1855
* NET  1124 = abc_11873_new_n1854
* NET  1125 = abc_11873_new_n1853
* NET  1126 = abc_11873_new_n1852
* NET  1127 = abc_11873_new_n1851
* NET  1128 = abc_11873_new_n1850
* NET  1129 = abc_11873_new_n1849
* NET  1130 = abc_11873_new_n1848
* NET  1131 = abc_11873_new_n1847
* NET  1132 = abc_11873_new_n1846
* NET  1133 = abc_11873_new_n1845
* NET  1134 = abc_11873_new_n1844
* NET  1135 = abc_11873_new_n1843
* NET  1136 = abc_11873_new_n1842
* NET  1137 = abc_11873_new_n1841
* NET  1138 = abc_11873_new_n1840
* NET  1139 = abc_11873_new_n1839
* NET  1140 = abc_11873_new_n1838
* NET  1141 = abc_11873_new_n1837
* NET  1142 = abc_11873_new_n1836
* NET  1143 = abc_11873_new_n1835
* NET  1144 = abc_11873_new_n1834
* NET  1145 = abc_11873_new_n1833
* NET  1146 = abc_11873_new_n1832
* NET  1147 = abc_11873_new_n1831
* NET  1148 = abc_11873_new_n1830
* NET  1149 = abc_11873_new_n1829
* NET  1150 = abc_11873_new_n1828
* NET  1151 = abc_11873_new_n1827
* NET  1152 = abc_11873_new_n1825
* NET  1153 = abc_11873_new_n1824
* NET  1154 = abc_11873_new_n1823
* NET  1155 = abc_11873_new_n1822
* NET  1156 = abc_11873_new_n1821
* NET  1157 = abc_11873_new_n1820
* NET  1158 = abc_11873_new_n1819
* NET  1159 = abc_11873_new_n1818
* NET  1160 = abc_11873_new_n1817
* NET  1161 = abc_11873_new_n1816
* NET  1162 = abc_11873_new_n1815
* NET  1163 = abc_11873_new_n1814
* NET  1164 = abc_11873_new_n1813
* NET  1165 = abc_11873_new_n1812
* NET  1166 = abc_11873_new_n1811
* NET  1167 = abc_11873_new_n1810
* NET  1168 = abc_11873_new_n1809
* NET  1169 = abc_11873_new_n1808
* NET  1170 = abc_11873_new_n1807
* NET  1171 = abc_11873_new_n1806
* NET  1172 = abc_11873_new_n1805
* NET  1173 = abc_11873_new_n1804
* NET  1174 = abc_11873_new_n1803
* NET  1175 = abc_11873_new_n1802
* NET  1176 = abc_11873_new_n1801
* NET  1177 = abc_11873_new_n1800
* NET  1178 = abc_11873_new_n1799
* NET  1179 = abc_11873_new_n1798
* NET  1180 = abc_11873_new_n1797
* NET  1181 = abc_11873_new_n1796
* NET  1182 = abc_11873_new_n1795
* NET  1183 = abc_11873_new_n1794
* NET  1184 = abc_11873_new_n1793
* NET  1185 = abc_11873_new_n1792
* NET  1186 = abc_11873_new_n1791
* NET  1187 = abc_11873_new_n1790
* NET  1188 = abc_11873_new_n1789
* NET  1189 = abc_11873_new_n1788
* NET  1190 = abc_11873_new_n1787
* NET  1191 = abc_11873_new_n1786
* NET  1192 = abc_11873_new_n1785
* NET  1193 = abc_11873_new_n1784
* NET  1194 = abc_11873_new_n1783
* NET  1195 = abc_11873_new_n1782
* NET  1196 = abc_11873_new_n1781
* NET  1197 = abc_11873_new_n1780
* NET  1198 = abc_11873_new_n1779
* NET  1199 = abc_11873_new_n1778
* NET  1200 = abc_11873_new_n1777
* NET  1201 = abc_11873_new_n1776
* NET  1202 = abc_11873_new_n1775
* NET  1203 = abc_11873_new_n1774
* NET  1204 = abc_11873_new_n1773
* NET  1205 = abc_11873_new_n1772
* NET  1206 = abc_11873_new_n1771
* NET  1207 = abc_11873_new_n1770
* NET  1208 = abc_11873_new_n1769
* NET  1209 = abc_11873_new_n1768
* NET  1210 = abc_11873_new_n1767
* NET  1211 = abc_11873_new_n1766
* NET  1212 = abc_11873_new_n1765
* NET  1213 = abc_11873_new_n1764
* NET  1214 = abc_11873_new_n1763
* NET  1215 = abc_11873_new_n1762
* NET  1216 = abc_11873_new_n1761
* NET  1217 = abc_11873_new_n1760
* NET  1218 = abc_11873_new_n1759
* NET  1219 = abc_11873_new_n1758
* NET  1220 = abc_11873_new_n1757
* NET  1221 = abc_11873_new_n1756
* NET  1222 = abc_11873_new_n1755
* NET  1223 = abc_11873_new_n1754
* NET  1224 = abc_11873_new_n1753
* NET  1225 = abc_11873_new_n1752
* NET  1226 = abc_11873_new_n1751
* NET  1227 = abc_11873_new_n1750
* NET  1228 = abc_11873_new_n1749
* NET  1229 = abc_11873_new_n1747
* NET  1230 = abc_11873_new_n1746
* NET  1231 = abc_11873_new_n1745
* NET  1232 = abc_11873_new_n1744
* NET  1233 = abc_11873_new_n1743
* NET  1234 = abc_11873_new_n1742
* NET  1235 = abc_11873_new_n1741
* NET  1236 = abc_11873_new_n1740
* NET  1237 = abc_11873_new_n1738
* NET  1238 = abc_11873_new_n1737
* NET  1239 = abc_11873_new_n1736
* NET  1240 = abc_11873_new_n1735
* NET  1241 = abc_11873_new_n1734
* NET  1242 = abc_11873_new_n1733
* NET  1243 = abc_11873_new_n1732
* NET  1244 = abc_11873_new_n1731
* NET  1245 = abc_11873_new_n1730
* NET  1246 = abc_11873_new_n1729
* NET  1247 = abc_11873_new_n1727
* NET  1248 = abc_11873_new_n1726
* NET  1249 = abc_11873_new_n1725
* NET  1250 = abc_11873_new_n1724
* NET  1251 = abc_11873_new_n1723
* NET  1252 = abc_11873_new_n1722
* NET  1253 = abc_11873_new_n1721
* NET  1254 = abc_11873_new_n1720
* NET  1255 = abc_11873_new_n1719
* NET  1256 = abc_11873_new_n1718
* NET  1257 = abc_11873_new_n1717
* NET  1258 = abc_11873_new_n1716
* NET  1259 = abc_11873_new_n1714
* NET  1260 = abc_11873_new_n1713
* NET  1261 = abc_11873_new_n1712
* NET  1262 = abc_11873_new_n1711
* NET  1263 = abc_11873_new_n1710
* NET  1264 = abc_11873_new_n1709
* NET  1265 = abc_11873_new_n1708
* NET  1266 = abc_11873_new_n1707
* NET  1267 = abc_11873_new_n1706
* NET  1268 = abc_11873_new_n1704
* NET  1269 = abc_11873_new_n1703
* NET  1270 = abc_11873_new_n1702
* NET  1271 = abc_11873_new_n1701
* NET  1272 = abc_11873_new_n1700
* NET  1273 = abc_11873_new_n1699
* NET  1274 = abc_11873_new_n1698
* NET  1275 = abc_11873_new_n1697
* NET  1276 = abc_11873_new_n1696
* NET  1277 = abc_11873_new_n1695
* NET  1278 = abc_11873_new_n1693
* NET  1279 = abc_11873_new_n1692
* NET  1280 = abc_11873_new_n1691
* NET  1281 = abc_11873_new_n1690
* NET  1282 = abc_11873_new_n1689
* NET  1283 = abc_11873_new_n1688
* NET  1284 = abc_11873_new_n1687
* NET  1285 = abc_11873_new_n1686
* NET  1286 = abc_11873_new_n1685
* NET  1287 = abc_11873_new_n1684
* NET  1288 = abc_11873_new_n1683
* NET  1289 = abc_11873_new_n1682
* NET  1290 = abc_11873_new_n1680
* NET  1291 = abc_11873_new_n1679
* NET  1292 = abc_11873_new_n1678
* NET  1293 = abc_11873_new_n1677
* NET  1294 = abc_11873_new_n1676
* NET  1295 = abc_11873_new_n1675
* NET  1296 = abc_11873_new_n1674
* NET  1297 = abc_11873_new_n1673
* NET  1298 = abc_11873_new_n1672
* NET  1299 = abc_11873_new_n1670
* NET  1300 = abc_11873_new_n1669
* NET  1301 = abc_11873_new_n1668
* NET  1302 = abc_11873_new_n1667
* NET  1303 = abc_11873_new_n1666
* NET  1304 = abc_11873_new_n1665
* NET  1305 = abc_11873_new_n1664
* NET  1306 = abc_11873_new_n1663
* NET  1307 = abc_11873_new_n1662
* NET  1308 = abc_11873_new_n1661
* NET  1309 = abc_11873_new_n1660
* NET  1310 = abc_11873_new_n1658
* NET  1311 = abc_11873_new_n1657
* NET  1312 = abc_11873_new_n1656
* NET  1313 = abc_11873_new_n1655
* NET  1314 = abc_11873_new_n1654
* NET  1315 = abc_11873_new_n1653
* NET  1316 = abc_11873_new_n1652
* NET  1317 = abc_11873_new_n1651
* NET  1318 = abc_11873_new_n1649
* NET  1319 = abc_11873_new_n1648
* NET  1320 = abc_11873_new_n1647
* NET  1321 = abc_11873_new_n1646
* NET  1322 = abc_11873_new_n1645
* NET  1323 = abc_11873_new_n1644
* NET  1324 = abc_11873_new_n1643
* NET  1325 = abc_11873_new_n1642
* NET  1326 = abc_11873_new_n1640
* NET  1327 = abc_11873_new_n1639
* NET  1328 = abc_11873_new_n1638
* NET  1329 = abc_11873_new_n1637
* NET  1330 = abc_11873_new_n1636
* NET  1331 = abc_11873_new_n1635
* NET  1332 = abc_11873_new_n1634
* NET  1333 = abc_11873_new_n1633
* NET  1334 = abc_11873_new_n1632
* NET  1335 = abc_11873_new_n1630
* NET  1336 = abc_11873_new_n1629
* NET  1337 = abc_11873_new_n1628
* NET  1338 = abc_11873_new_n1627
* NET  1339 = abc_11873_new_n1626
* NET  1340 = abc_11873_new_n1625
* NET  1341 = abc_11873_new_n1624
* NET  1342 = abc_11873_new_n1623
* NET  1343 = abc_11873_new_n1622
* NET  1344 = abc_11873_new_n1620
* NET  1345 = abc_11873_new_n1619
* NET  1346 = abc_11873_new_n1618
* NET  1347 = abc_11873_new_n1617
* NET  1348 = abc_11873_new_n1616
* NET  1349 = abc_11873_new_n1615
* NET  1350 = abc_11873_new_n1614
* NET  1351 = abc_11873_new_n1613
* NET  1352 = abc_11873_new_n1611
* NET  1353 = abc_11873_new_n1610
* NET  1354 = abc_11873_new_n1609
* NET  1355 = abc_11873_new_n1608
* NET  1356 = abc_11873_new_n1607
* NET  1357 = abc_11873_new_n1606
* NET  1358 = abc_11873_new_n1605
* NET  1359 = abc_11873_new_n1604
* NET  1360 = abc_11873_new_n1603
* NET  1361 = abc_11873_new_n1602
* NET  1362 = abc_11873_new_n1601
* NET  1363 = abc_11873_new_n1599
* NET  1364 = abc_11873_new_n1598
* NET  1365 = abc_11873_new_n1597
* NET  1366 = abc_11873_new_n1596
* NET  1367 = abc_11873_new_n1595
* NET  1368 = abc_11873_new_n1594
* NET  1369 = abc_11873_new_n1593
* NET  1370 = abc_11873_new_n1592
* NET  1371 = abc_11873_new_n1590
* NET  1372 = abc_11873_new_n1589
* NET  1373 = abc_11873_new_n1588
* NET  1374 = abc_11873_new_n1587
* NET  1375 = abc_11873_new_n1586
* NET  1376 = abc_11873_new_n1585
* NET  1377 = abc_11873_new_n1584
* NET  1378 = abc_11873_new_n1583
* NET  1379 = abc_11873_new_n1582
* NET  1380 = abc_11873_new_n1581
* NET  1381 = abc_11873_new_n1580
* NET  1382 = abc_11873_new_n1579
* NET  1383 = abc_11873_new_n1578
* NET  1384 = abc_11873_new_n1577
* NET  1385 = abc_11873_new_n1576
* NET  1386 = abc_11873_new_n1575
* NET  1387 = abc_11873_new_n1574
* NET  1388 = abc_11873_new_n1573
* NET  1389 = abc_11873_new_n1572
* NET  1390 = abc_11873_new_n1571
* NET  1391 = abc_11873_new_n1570
* NET  1392 = abc_11873_new_n1569
* NET  1393 = abc_11873_new_n1568
* NET  1394 = abc_11873_new_n1551
* NET  1395 = abc_11873_new_n1550
* NET  1396 = abc_11873_new_n1549
* NET  1397 = abc_11873_new_n1548
* NET  1398 = abc_11873_new_n1547
* NET  1399 = abc_11873_new_n1546
* NET  1400 = abc_11873_new_n1545
* NET  1401 = abc_11873_new_n1544
* NET  1402 = abc_11873_new_n1543
* NET  1403 = abc_11873_new_n1542
* NET  1404 = abc_11873_new_n1541
* NET  1405 = abc_11873_new_n1540
* NET  1406 = abc_11873_new_n1539
* NET  1407 = abc_11873_new_n1538
* NET  1408 = abc_11873_new_n1537
* NET  1409 = abc_11873_new_n1536
* NET  1410 = abc_11873_new_n1535
* NET  1411 = abc_11873_new_n1534
* NET  1412 = abc_11873_new_n1533
* NET  1413 = abc_11873_new_n1532
* NET  1414 = abc_11873_new_n1531
* NET  1415 = abc_11873_new_n1530
* NET  1416 = abc_11873_new_n1529
* NET  1417 = abc_11873_new_n1528
* NET  1418 = abc_11873_new_n1527
* NET  1419 = abc_11873_new_n1526
* NET  1420 = abc_11873_new_n1525
* NET  1421 = abc_11873_new_n1524
* NET  1422 = abc_11873_new_n1523
* NET  1423 = abc_11873_new_n1522
* NET  1424 = abc_11873_new_n1521
* NET  1425 = abc_11873_new_n1520
* NET  1426 = abc_11873_new_n1519
* NET  1427 = abc_11873_new_n1518
* NET  1428 = abc_11873_new_n1517
* NET  1429 = abc_11873_new_n1516
* NET  1430 = abc_11873_new_n1515
* NET  1431 = abc_11873_new_n1514
* NET  1432 = abc_11873_new_n1513
* NET  1433 = abc_11873_new_n1512
* NET  1434 = abc_11873_new_n1511
* NET  1435 = abc_11873_new_n1510
* NET  1436 = abc_11873_new_n1509
* NET  1437 = abc_11873_new_n1508
* NET  1438 = abc_11873_new_n1507
* NET  1439 = abc_11873_new_n1506
* NET  1440 = abc_11873_new_n1505
* NET  1441 = abc_11873_new_n1504
* NET  1442 = abc_11873_new_n1503
* NET  1443 = abc_11873_new_n1502
* NET  1444 = abc_11873_new_n1499
* NET  1445 = abc_11873_new_n1498
* NET  1446 = abc_11873_new_n1497
* NET  1447 = abc_11873_new_n1496
* NET  1448 = abc_11873_new_n1495
* NET  1449 = abc_11873_new_n1494
* NET  1450 = abc_11873_new_n1493
* NET  1451 = abc_11873_new_n1492
* NET  1452 = abc_11873_new_n1491
* NET  1453 = abc_11873_new_n1489
* NET  1454 = abc_11873_new_n1488
* NET  1455 = abc_11873_new_n1487
* NET  1456 = abc_11873_new_n1486
* NET  1457 = abc_11873_new_n1485
* NET  1458 = abc_11873_new_n1484
* NET  1459 = abc_11873_new_n1483
* NET  1460 = abc_11873_new_n1482
* NET  1461 = abc_11873_new_n1481
* NET  1462 = abc_11873_new_n1479
* NET  1463 = abc_11873_new_n1478
* NET  1464 = abc_11873_new_n1477
* NET  1465 = abc_11873_new_n1476
* NET  1466 = abc_11873_new_n1475
* NET  1467 = abc_11873_new_n1474
* NET  1468 = abc_11873_new_n1473
* NET  1469 = abc_11873_new_n1471
* NET  1470 = abc_11873_new_n1470
* NET  1471 = abc_11873_new_n1469
* NET  1472 = abc_11873_new_n1468
* NET  1473 = abc_11873_new_n1466
* NET  1474 = abc_11873_new_n1465
* NET  1475 = abc_11873_new_n1464
* NET  1476 = abc_11873_new_n1463
* NET  1477 = abc_11873_new_n1462
* NET  1478 = abc_11873_new_n1461
* NET  1479 = abc_11873_new_n1460
* NET  1480 = abc_11873_new_n1459
* NET  1481 = abc_11873_new_n1457
* NET  1482 = abc_11873_new_n1456
* NET  1483 = abc_11873_new_n1455
* NET  1484 = abc_11873_new_n1454
* NET  1485 = abc_11873_new_n1453
* NET  1486 = abc_11873_new_n1452
* NET  1487 = abc_11873_new_n1451
* NET  1488 = abc_11873_new_n1450
* NET  1489 = abc_11873_new_n1449
* NET  1490 = abc_11873_new_n1448
* NET  1491 = abc_11873_new_n1447
* NET  1492 = abc_11873_new_n1446
* NET  1493 = abc_11873_new_n1436
* NET  1494 = abc_11873_new_n1435
* NET  1495 = abc_11873_new_n1434
* NET  1496 = abc_11873_new_n1432
* NET  1497 = abc_11873_new_n1431
* NET  1498 = abc_11873_new_n1430
* NET  1499 = abc_11873_new_n1429
* NET  1500 = abc_11873_new_n1428
* NET  1501 = abc_11873_new_n1427
* NET  1502 = abc_11873_new_n1426
* NET  1503 = abc_11873_new_n1425
* NET  1504 = abc_11873_new_n1424
* NET  1505 = abc_11873_new_n1423
* NET  1506 = abc_11873_new_n1420
* NET  1507 = abc_11873_new_n1419
* NET  1508 = abc_11873_new_n1418
* NET  1509 = abc_11873_new_n1417
* NET  1510 = abc_11873_new_n1416
* NET  1511 = abc_11873_new_n1414
* NET  1512 = abc_11873_new_n1413
* NET  1513 = abc_11873_new_n1412
* NET  1514 = abc_11873_new_n1411
* NET  1515 = abc_11873_new_n1410
* NET  1516 = abc_11873_new_n1409
* NET  1517 = abc_11873_new_n1407
* NET  1518 = abc_11873_new_n1406
* NET  1519 = abc_11873_new_n1405
* NET  1520 = abc_11873_new_n1404
* NET  1521 = abc_11873_new_n1403
* NET  1522 = abc_11873_new_n1402
* NET  1523 = abc_11873_new_n1401
* NET  1524 = abc_11873_new_n1399
* NET  1525 = abc_11873_new_n1398
* NET  1526 = abc_11873_new_n1397
* NET  1527 = abc_11873_new_n1396
* NET  1528 = abc_11873_new_n1395
* NET  1529 = abc_11873_new_n1394
* NET  1530 = abc_11873_new_n1393
* NET  1531 = abc_11873_new_n1392
* NET  1532 = abc_11873_new_n1391
* NET  1533 = abc_11873_new_n1390
* NET  1534 = abc_11873_new_n1388
* NET  1535 = abc_11873_new_n1387
* NET  1536 = abc_11873_new_n1386
* NET  1537 = abc_11873_new_n1384
* NET  1538 = abc_11873_new_n1383
* NET  1539 = abc_11873_new_n1382
* NET  1540 = abc_11873_new_n1380
* NET  1541 = abc_11873_new_n1378
* NET  1542 = abc_11873_new_n1376
* NET  1543 = abc_11873_new_n1375
* NET  1544 = abc_11873_new_n1374
* NET  1545 = abc_11873_new_n1373
* NET  1546 = abc_11873_new_n1372
* NET  1547 = abc_11873_new_n1369
* NET  1548 = abc_11873_new_n1367
* NET  1549 = abc_11873_new_n1366
* NET  1550 = abc_11873_new_n1365
* NET  1551 = abc_11873_new_n1364
* NET  1552 = abc_11873_new_n1363
* NET  1553 = abc_11873_new_n1362
* NET  1554 = abc_11873_new_n1361
* NET  1555 = abc_11873_new_n1359
* NET  1556 = abc_11873_new_n1358
* NET  1557 = abc_11873_new_n1357
* NET  1558 = abc_11873_new_n1354
* NET  1559 = abc_11873_new_n1353
* NET  1560 = abc_11873_new_n1352
* NET  1561 = abc_11873_new_n1351
* NET  1562 = abc_11873_new_n1350
* NET  1563 = abc_11873_new_n1347
* NET  1564 = abc_11873_new_n1345
* NET  1565 = abc_11873_new_n1344
* NET  1566 = abc_11873_new_n1343
* NET  1567 = abc_11873_new_n1342
* NET  1568 = abc_11873_new_n1341
* NET  1569 = abc_11873_new_n1339
* NET  1570 = abc_11873_new_n1338
* NET  1571 = abc_11873_new_n1337
* NET  1572 = abc_11873_new_n1336
* NET  1573 = abc_11873_new_n1335
* NET  1574 = abc_11873_new_n1334
* NET  1575 = abc_11873_new_n1333
* NET  1576 = abc_11873_new_n1332
* NET  1577 = abc_11873_new_n1331
* NET  1578 = abc_11873_new_n1330
* NET  1579 = abc_11873_new_n1329
* NET  1580 = abc_11873_new_n1328
* NET  1581 = abc_11873_new_n1327
* NET  1582 = abc_11873_new_n1326
* NET  1583 = abc_11873_new_n1325
* NET  1584 = abc_11873_new_n1324
* NET  1585 = abc_11873_new_n1323
* NET  1586 = abc_11873_new_n1322
* NET  1587 = abc_11873_new_n1321
* NET  1588 = abc_11873_new_n1320
* NET  1589 = abc_11873_new_n1319
* NET  1590 = abc_11873_new_n1318
* NET  1591 = abc_11873_new_n1317
* NET  1592 = abc_11873_new_n1316
* NET  1593 = abc_11873_new_n1315
* NET  1594 = abc_11873_new_n1314
* NET  1595 = abc_11873_new_n1313
* NET  1596 = abc_11873_new_n1311
* NET  1597 = abc_11873_new_n1310
* NET  1598 = abc_11873_new_n1308
* NET  1599 = abc_11873_new_n1307
* NET  1600 = abc_11873_new_n1306
* NET  1601 = abc_11873_new_n1305
* NET  1602 = abc_11873_new_n1303
* NET  1603 = abc_11873_new_n1302
* NET  1604 = abc_11873_new_n1300
* NET  1605 = abc_11873_new_n1299
* NET  1606 = abc_11873_new_n1297
* NET  1607 = abc_11873_new_n1296
* NET  1608 = abc_11873_new_n1294
* NET  1609 = abc_11873_new_n1293
* NET  1610 = abc_11873_new_n1292
* NET  1611 = abc_11873_new_n1290
* NET  1612 = abc_11873_new_n1289
* NET  1613 = abc_11873_new_n1287
* NET  1614 = abc_11873_new_n1286
* NET  1615 = abc_11873_new_n1285
* NET  1616 = abc_11873_new_n1283
* NET  1617 = abc_11873_new_n1282
* NET  1618 = abc_11873_new_n1280
* NET  1619 = abc_11873_new_n1279
* NET  1620 = abc_11873_new_n1278
* NET  1621 = abc_11873_new_n1273
* NET  1622 = abc_11873_new_n1264
* NET  1623 = abc_11873_new_n1255
* NET  1624 = abc_11873_new_n1246
* NET  1625 = abc_11873_new_n1244
* NET  1626 = abc_11873_new_n1243
* NET  1627 = abc_11873_new_n1242
* NET  1628 = abc_11873_new_n1241
* NET  1629 = abc_11873_new_n1239
* NET  1630 = abc_11873_new_n1238
* NET  1631 = abc_11873_new_n1237
* NET  1632 = abc_11873_new_n1236
* NET  1633 = abc_11873_new_n1235
* NET  1634 = abc_11873_new_n1233
* NET  1635 = abc_11873_new_n1232
* NET  1636 = abc_11873_new_n1231
* NET  1637 = abc_11873_new_n1230
* NET  1638 = abc_11873_new_n1229
* NET  1639 = abc_11873_new_n1228
* NET  1640 = abc_11873_new_n1227
* NET  1641 = abc_11873_new_n1226
* NET  1642 = abc_11873_new_n1224
* NET  1643 = abc_11873_new_n1222
* NET  1644 = abc_11873_new_n1221
* NET  1645 = abc_11873_new_n1220
* NET  1646 = abc_11873_new_n1219
* NET  1647 = abc_11873_new_n1217
* NET  1648 = abc_11873_new_n1216
* NET  1649 = abc_11873_new_n1215
* NET  1650 = abc_11873_new_n1214
* NET  1651 = abc_11873_new_n1213
* NET  1652 = abc_11873_new_n1211
* NET  1653 = abc_11873_new_n1210
* NET  1654 = abc_11873_new_n1209
* NET  1655 = abc_11873_new_n1208
* NET  1656 = abc_11873_new_n1207
* NET  1657 = abc_11873_new_n1206
* NET  1658 = abc_11873_new_n1205
* NET  1659 = abc_11873_new_n1204
* NET  1660 = abc_11873_new_n1203
* NET  1661 = abc_11873_new_n1201
* NET  1662 = abc_11873_new_n1200
* NET  1663 = abc_11873_new_n1199
* NET  1664 = abc_11873_new_n1198
* NET  1665 = abc_11873_new_n1197
* NET  1666 = abc_11873_new_n1196
* NET  1667 = abc_11873_new_n1195
* NET  1668 = abc_11873_new_n1194
* NET  1669 = abc_11873_new_n1191
* NET  1670 = abc_11873_new_n1190
* NET  1671 = abc_11873_new_n1189
* NET  1672 = abc_11873_new_n1188
* NET  1673 = abc_11873_new_n1187
* NET  1674 = abc_11873_new_n1185
* NET  1675 = abc_11873_new_n1184
* NET  1676 = abc_11873_new_n1183
* NET  1677 = abc_11873_new_n1182
* NET  1678 = abc_11873_new_n1181
* NET  1679 = abc_11873_new_n1179
* NET  1680 = abc_11873_new_n1178
* NET  1681 = abc_11873_new_n1177
* NET  1682 = abc_11873_new_n1176
* NET  1683 = abc_11873_new_n1175
* NET  1684 = abc_11873_new_n1173
* NET  1685 = abc_11873_new_n1172
* NET  1686 = abc_11873_new_n1171
* NET  1687 = abc_11873_new_n1170
* NET  1688 = abc_11873_new_n1169
* NET  1689 = abc_11873_new_n1167
* NET  1690 = abc_11873_new_n1166
* NET  1691 = abc_11873_new_n1165
* NET  1692 = abc_11873_new_n1164
* NET  1693 = abc_11873_new_n1163
* NET  1694 = abc_11873_new_n1161
* NET  1695 = abc_11873_new_n1160
* NET  1696 = abc_11873_new_n1159
* NET  1697 = abc_11873_new_n1158
* NET  1698 = abc_11873_new_n1157
* NET  1699 = abc_11873_new_n1155
* NET  1700 = abc_11873_new_n1154
* NET  1701 = abc_11873_new_n1153
* NET  1702 = abc_11873_new_n1152
* NET  1703 = abc_11873_new_n1151
* NET  1704 = abc_11873_new_n1149
* NET  1705 = abc_11873_new_n1148
* NET  1706 = abc_11873_new_n1147
* NET  1707 = abc_11873_new_n1146
* NET  1708 = abc_11873_new_n1145
* NET  1709 = abc_11873_new_n1144
* NET  1710 = abc_11873_new_n1142
* NET  1711 = abc_11873_new_n1141
* NET  1712 = abc_11873_new_n1140
* NET  1713 = abc_11873_new_n1139
* NET  1714 = abc_11873_new_n1138
* NET  1715 = abc_11873_new_n1137
* NET  1716 = abc_11873_new_n1136
* NET  1717 = abc_11873_new_n1134
* NET  1718 = abc_11873_new_n1133
* NET  1719 = abc_11873_new_n1132
* NET  1720 = abc_11873_new_n1131
* NET  1721 = abc_11873_new_n1130
* NET  1722 = abc_11873_new_n1129
* NET  1723 = abc_11873_new_n1128
* NET  1724 = abc_11873_new_n1126
* NET  1725 = abc_11873_new_n1125
* NET  1726 = abc_11873_new_n1124
* NET  1727 = abc_11873_new_n1123
* NET  1728 = abc_11873_new_n1122
* NET  1729 = abc_11873_new_n1121
* NET  1730 = abc_11873_new_n1120
* NET  1731 = abc_11873_new_n1119
* NET  1732 = abc_11873_new_n1117
* NET  1733 = abc_11873_new_n1116
* NET  1734 = abc_11873_new_n1115
* NET  1735 = abc_11873_new_n1114
* NET  1736 = abc_11873_new_n1113
* NET  1737 = abc_11873_new_n1112
* NET  1738 = abc_11873_new_n1111
* NET  1739 = abc_11873_new_n1109
* NET  1740 = abc_11873_new_n1108
* NET  1741 = abc_11873_new_n1107
* NET  1742 = abc_11873_new_n1106
* NET  1743 = abc_11873_new_n1105
* NET  1744 = abc_11873_new_n1104
* NET  1745 = abc_11873_new_n1103
* NET  1746 = abc_11873_new_n1101
* NET  1747 = abc_11873_new_n1100
* NET  1748 = abc_11873_new_n1099
* NET  1749 = abc_11873_new_n1098
* NET  1750 = abc_11873_new_n1097
* NET  1751 = abc_11873_new_n1096
* NET  1752 = abc_11873_new_n1095
* NET  1753 = abc_11873_new_n1093
* NET  1754 = abc_11873_new_n1092
* NET  1755 = abc_11873_new_n1091
* NET  1756 = abc_11873_new_n1090
* NET  1757 = abc_11873_new_n1089
* NET  1758 = abc_11873_new_n1088
* NET  1759 = abc_11873_new_n1087
* NET  1760 = abc_11873_new_n1085
* NET  1761 = abc_11873_new_n1084
* NET  1762 = abc_11873_new_n1083
* NET  1763 = abc_11873_new_n1082
* NET  1764 = abc_11873_new_n1081
* NET  1765 = abc_11873_new_n1080
* NET  1766 = abc_11873_new_n1079
* NET  1767 = abc_11873_new_n1078
* NET  1768 = abc_11873_new_n1077
* NET  1769 = abc_11873_new_n1076
* NET  1770 = abc_11873_new_n1075
* NET  1771 = abc_11873_new_n1074
* NET  1772 = abc_11873_new_n1073
* NET  1773 = abc_11873_new_n1072
* NET  1774 = abc_11873_new_n1071
* NET  1775 = abc_11873_new_n1070
* NET  1776 = abc_11873_new_n1069
* NET  1777 = abc_11873_new_n1068
* NET  1778 = abc_11873_new_n1067
* NET  1779 = abc_11873_new_n1066
* NET  1780 = abc_11873_new_n1065
* NET  1781 = abc_11873_new_n1064
* NET  1782 = abc_11873_new_n1063
* NET  1783 = abc_11873_new_n1062
* NET  1784 = abc_11873_new_n1061
* NET  1785 = abc_11873_new_n1060
* NET  1786 = abc_11873_new_n1059
* NET  1787 = abc_11873_new_n1058
* NET  1788 = abc_11873_new_n1057
* NET  1789 = abc_11873_new_n1056
* NET  1790 = abc_11873_new_n1055
* NET  1791 = abc_11873_new_n1054
* NET  1792 = abc_11873_new_n1053
* NET  1793 = abc_11873_new_n1052
* NET  1794 = abc_11873_new_n1050
* NET  1795 = abc_11873_new_n1049
* NET  1796 = abc_11873_new_n1048
* NET  1797 = abc_11873_new_n1047
* NET  1798 = abc_11873_new_n1046
* NET  1799 = abc_11873_new_n1045
* NET  1800 = abc_11873_new_n1044
* NET  1801 = abc_11873_new_n1043
* NET  1802 = abc_11873_new_n1042
* NET  1803 = abc_11873_new_n1041
* NET  1804 = abc_11873_new_n1040
* NET  1805 = abc_11873_new_n1038
* NET  1806 = abc_11873_new_n1037
* NET  1807 = abc_11873_new_n1036
* NET  1808 = abc_11873_new_n1035
* NET  1809 = abc_11873_new_n1034
* NET  1810 = abc_11873_new_n1033
* NET  1811 = abc_11873_new_n1032
* NET  1812 = abc_11873_new_n1031
* NET  1813 = abc_11873_new_n1030
* NET  1814 = abc_11873_new_n1029
* NET  1815 = abc_11873_new_n1028
* NET  1816 = abc_11873_new_n1026
* NET  1817 = abc_11873_new_n1025
* NET  1818 = abc_11873_new_n1024
* NET  1819 = abc_11873_new_n1023
* NET  1820 = abc_11873_new_n1022
* NET  1821 = abc_11873_new_n1021
* NET  1822 = abc_11873_new_n1020
* NET  1823 = abc_11873_new_n1019
* NET  1824 = abc_11873_new_n1018
* NET  1825 = abc_11873_new_n1017
* NET  1826 = abc_11873_new_n1016
* NET  1827 = abc_11873_new_n1015
* NET  1828 = abc_11873_new_n1013
* NET  1829 = abc_11873_new_n1012
* NET  1830 = abc_11873_new_n1011
* NET  1831 = abc_11873_new_n1010
* NET  1832 = abc_11873_new_n1009
* NET  1833 = abc_11873_new_n1008
* NET  1834 = abc_11873_new_n1007
* NET  1835 = abc_11873_new_n1006
* NET  1836 = abc_11873_new_n1005
* NET  1837 = abc_11873_new_n1004
* NET  1838 = abc_11873_new_n1003
* NET  1839 = abc_11873_new_n1001
* NET  1840 = abc_11873_new_n1000
* NET  1841 = abc_11873_flatten_mos6502_0_adj_bcd_0_0
* NET  1842 = abc_11873_auto_rtlil_cc_2560_muxgate_11872
* NET  1843 = abc_11873_auto_rtlil_cc_2560_muxgate_11870
* NET  1844 = abc_11873_auto_rtlil_cc_2560_muxgate_11868
* NET  1845 = abc_11873_auto_rtlil_cc_2560_muxgate_11866
* NET  1846 = abc_11873_auto_rtlil_cc_2560_muxgate_11864
* NET  1847 = abc_11873_auto_rtlil_cc_2560_muxgate_11862
* NET  1848 = abc_11873_auto_rtlil_cc_2560_muxgate_11860
* NET  1849 = abc_11873_auto_rtlil_cc_2560_muxgate_11858
* NET  1850 = abc_11873_auto_rtlil_cc_2560_muxgate_11856
* NET  1851 = abc_11873_auto_rtlil_cc_2560_muxgate_11854
* NET  1852 = abc_11873_auto_rtlil_cc_2560_muxgate_11852
* NET  1853 = abc_11873_auto_rtlil_cc_2560_muxgate_11850
* NET  1854 = abc_11873_auto_rtlil_cc_2560_muxgate_11848
* NET  1855 = abc_11873_auto_rtlil_cc_2560_muxgate_11846
* NET  1856 = abc_11873_auto_rtlil_cc_2560_muxgate_11844
* NET  1857 = abc_11873_auto_rtlil_cc_2560_muxgate_11842
* NET  1858 = abc_11873_auto_rtlil_cc_2560_muxgate_11840
* NET  1859 = abc_11873_auto_rtlil_cc_2560_muxgate_11838
* NET  1860 = abc_11873_auto_rtlil_cc_2560_muxgate_11836
* NET  1861 = abc_11873_auto_rtlil_cc_2560_muxgate_11834
* NET  1862 = abc_11873_auto_rtlil_cc_2560_muxgate_11832
* NET  1863 = abc_11873_auto_rtlil_cc_2560_muxgate_11830
* NET  1864 = abc_11873_auto_rtlil_cc_2560_muxgate_11828
* NET  1865 = abc_11873_auto_rtlil_cc_2560_muxgate_11826
* NET  1866 = abc_11873_auto_rtlil_cc_2560_muxgate_11824
* NET  1867 = abc_11873_auto_rtlil_cc_2560_muxgate_11822
* NET  1868 = abc_11873_auto_rtlil_cc_2560_muxgate_11820
* NET  1869 = abc_11873_auto_rtlil_cc_2560_muxgate_11818
* NET  1870 = abc_11873_auto_rtlil_cc_2560_muxgate_11816
* NET  1871 = abc_11873_auto_rtlil_cc_2560_muxgate_11814
* NET  1872 = abc_11873_auto_rtlil_cc_2560_muxgate_11812
* NET  1873 = abc_11873_auto_rtlil_cc_2560_muxgate_11810
* NET  1874 = abc_11873_auto_rtlil_cc_2560_muxgate_11808
* NET  1875 = abc_11873_auto_rtlil_cc_2560_muxgate_11806
* NET  1876 = abc_11873_auto_rtlil_cc_2560_muxgate_11804
* NET  1877 = abc_11873_auto_rtlil_cc_2560_muxgate_11802
* NET  1878 = abc_11873_auto_rtlil_cc_2560_muxgate_11800
* NET  1879 = abc_11873_auto_rtlil_cc_2560_muxgate_11798
* NET  1880 = abc_11873_auto_rtlil_cc_2560_muxgate_11796
* NET  1881 = abc_11873_auto_rtlil_cc_2560_muxgate_11794
* NET  1882 = abc_11873_auto_rtlil_cc_2560_muxgate_11792
* NET  1883 = abc_11873_auto_rtlil_cc_2560_muxgate_11790
* NET  1884 = abc_11873_auto_rtlil_cc_2560_muxgate_11788
* NET  1885 = abc_11873_auto_rtlil_cc_2560_muxgate_11786
* NET  1886 = abc_11873_auto_rtlil_cc_2560_muxgate_11784
* NET  1887 = abc_11873_auto_rtlil_cc_2560_muxgate_11782
* NET  1888 = abc_11873_auto_rtlil_cc_2560_muxgate_11780
* NET  1889 = abc_11873_auto_rtlil_cc_2560_muxgate_11778
* NET  1890 = abc_11873_auto_rtlil_cc_2560_muxgate_11776
* NET  1891 = abc_11873_auto_rtlil_cc_2560_muxgate_11774
* NET  1892 = abc_11873_auto_rtlil_cc_2560_muxgate_11770
* NET  1893 = abc_11873_auto_rtlil_cc_2560_muxgate_11768
* NET  1894 = abc_11873_auto_rtlil_cc_2560_muxgate_11766
* NET  1895 = abc_11873_auto_rtlil_cc_2560_muxgate_11764
* NET  1896 = abc_11873_auto_rtlil_cc_2560_muxgate_11762
* NET  1897 = abc_11873_auto_rtlil_cc_2560_muxgate_11760
* NET  1898 = abc_11873_auto_rtlil_cc_2560_muxgate_11758
* NET  1899 = abc_11873_auto_rtlil_cc_2560_muxgate_11756
* NET  1900 = abc_11873_auto_rtlil_cc_2560_muxgate_11754
* NET  1901 = abc_11873_auto_rtlil_cc_2560_muxgate_11752
* NET  1902 = abc_11873_auto_rtlil_cc_2560_muxgate_11748
* NET  1903 = abc_11873_auto_rtlil_cc_2560_muxgate_11746
* NET  1904 = abc_11873_auto_rtlil_cc_2560_muxgate_11742
* NET  1905 = abc_11873_auto_rtlil_cc_2560_muxgate_11740
* NET  1906 = abc_11873_auto_rtlil_cc_2560_muxgate_11738
* NET  1907 = abc_11873_auto_rtlil_cc_2560_muxgate_11736
* NET  1908 = abc_11873_auto_rtlil_cc_2560_muxgate_11734
* NET  1909 = abc_11873_auto_rtlil_cc_2560_muxgate_11732
* NET  1910 = abc_11873_auto_rtlil_cc_2560_muxgate_11730
* NET  1911 = abc_11873_auto_rtlil_cc_2560_muxgate_11728
* NET  1912 = abc_11873_auto_rtlil_cc_2560_muxgate_11726
* NET  1913 = abc_11873_auto_rtlil_cc_2560_muxgate_11724
* NET  1914 = abc_11873_auto_rtlil_cc_2560_muxgate_11722
* NET  1915 = abc_11873_auto_rtlil_cc_2560_muxgate_11720
* NET  1916 = abc_11873_auto_rtlil_cc_2560_muxgate_11716
* NET  1917 = abc_11873_auto_rtlil_cc_2560_muxgate_11714
* NET  1918 = abc_11873_auto_rtlil_cc_2560_muxgate_11712
* NET  1919 = abc_11873_auto_rtlil_cc_2560_muxgate_11710
* NET  1920 = abc_11873_auto_rtlil_cc_2560_muxgate_11708
* NET  1921 = abc_11873_auto_rtlil_cc_2560_muxgate_11706
* NET  1922 = abc_11873_auto_rtlil_cc_2560_muxgate_11704
* NET  1923 = abc_11873_auto_rtlil_cc_2560_muxgate_11702
* NET  1924 = abc_11873_auto_rtlil_cc_2560_muxgate_11700
* NET  1925 = abc_11873_auto_rtlil_cc_2560_muxgate_11698
* NET  1926 = abc_11873_auto_rtlil_cc_2560_muxgate_11696
* NET  1927 = abc_11873_auto_rtlil_cc_2560_muxgate_11694
* NET  1928 = abc_11873_auto_rtlil_cc_2560_muxgate_11692
* NET  1929 = abc_11873_auto_rtlil_cc_2560_muxgate_11690
* NET  1930 = abc_11873_auto_rtlil_cc_2560_muxgate_11688
* NET  1931 = abc_11873_auto_rtlil_cc_2560_muxgate_11686
* NET  1932 = abc_11873_auto_rtlil_cc_2560_muxgate_11684
* NET  1933 = abc_11873_auto_rtlil_cc_2560_muxgate_11682
* NET  1934 = abc_11873_auto_rtlil_cc_2560_muxgate_11680
* NET  1935 = abc_11873_auto_rtlil_cc_2560_muxgate_11678
* NET  1936 = abc_11873_auto_rtlil_cc_2560_muxgate_11676
* NET  1937 = abc_11873_auto_rtlil_cc_2560_muxgate_11672
* NET  1938 = abc_11873_auto_rtlil_cc_2560_muxgate_11670
* NET  1939 = abc_11873_auto_rtlil_cc_2560_muxgate_11668
* NET  1940 = abc_11873_auto_rtlil_cc_2560_muxgate_11666
* NET  1941 = abc_11873_auto_rtlil_cc_2560_muxgate_11664
* NET  1942 = abc_11873_auto_rtlil_cc_2560_muxgate_11662
* NET  1943 = abc_11873_auto_rtlil_cc_2560_muxgate_11660
* NET  1944 = abc_11873_auto_rtlil_cc_2560_muxgate_11658
* NET  1945 = abc_11873_auto_rtlil_cc_2560_muxgate_11656
* NET  1946 = abc_11873_auto_rtlil_cc_2560_muxgate_11654
* NET  1947 = abc_11873_auto_rtlil_cc_2560_muxgate_11652
* NET  1948 = abc_11873_auto_rtlil_cc_2560_muxgate_11650
* NET  1949 = abc_11873_auto_rtlil_cc_2560_muxgate_11648
* NET  1950 = abc_11873_auto_rtlil_cc_2560_muxgate_11646
* NET  1951 = abc_11873_auto_rtlil_cc_2560_muxgate_11644
* NET  1952 = abc_11873_auto_rtlil_cc_2560_muxgate_11642
* NET  1953 = abc_11873_auto_rtlil_cc_2560_muxgate_11640
* NET  1954 = abc_11873_auto_rtlil_cc_2560_muxgate_11638
* NET  1955 = abc_11873_auto_rtlil_cc_2560_muxgate_11636
* NET  1956 = abc_11873_auto_rtlil_cc_2560_muxgate_11634
* NET  1957 = abc_11873_auto_rtlil_cc_2560_muxgate_11632
* NET  1958 = abc_11873_auto_rtlil_cc_2560_muxgate_11630
* NET  1959 = abc_11873_auto_rtlil_cc_2560_muxgate_11628
* NET  1960 = abc_11873_auto_rtlil_cc_2560_muxgate_11626
* NET  1961 = abc_11873_auto_rtlil_cc_2560_muxgate_11624
* NET  1962 = abc_11873_auto_rtlil_cc_2560_muxgate_11622
* NET  1963 = abc_11873_auto_rtlil_cc_2560_muxgate_11620
* NET  1964 = abc_11873_auto_rtlil_cc_2560_muxgate_11618
* NET  1965 = abc_11873_auto_rtlil_cc_2560_muxgate_11616
* NET  1966 = abc_11873_auto_rtlil_cc_2560_muxgate_11614
* NET  1967 = abc_11873_auto_rtlil_cc_2560_muxgate_11612
* NET  1968 = abc_11873_auto_rtlil_cc_2560_muxgate_11610
* NET  1969 = a[9]
* NET  1970 = a[8]
* NET  1971 = a[7]
* NET  1972 = a[6]
* NET  1973 = a[5]
* NET  1974 = a[4]
* NET  1975 = a[3]
* NET  1976 = a[2]
* NET  1977 = a[15]
* NET  1978 = a[14]
* NET  1979 = a[13]
* NET  1980 = a[12]
* NET  1981 = a[11]
* NET  1982 = a[10]
* NET  1983 = a[1]
* NET  1984 = a[0]

xfeed_369 2 1 decap_w0
xfeed_368 2 1 decap_w0
xfeed_367 2 1 decap_w0
xfeed_366 2 1 decap_w0
xfeed_365 2 1 decap_w0
xfeed_364 2 1 decap_w0
xfeed_363 2 1 decap_w0
xfeed_362 2 1 decap_w0
xfeed_361 2 1 decap_w0
xfeed_360 2 1 decap_w0
xsubckt_458_o2_x2 1 424 2 525 677 o2_x2
xsubckt_463_mx2_x2 1 419 2 103 13 11 mx2_x2
xsubckt_464_mx2_x2 1 418 2 103 66 111 mx2_x2
xsubckt_465_mx2_x2 1 417 2 104 418 419 mx2_x2
xsubckt_495_ao22_x2 1 388 2 755 760 780 ao22_x2
xsubckt_1285_a3_x2 2 1355 1 1356 1364 1373 a3_x2
xsubckt_1450_a3_x2 2 1204 1 530 568 585 a3_x2
xsubckt_1461_oa22_x2 1 1193 2 1799 1205 1195 oa22_x2
xsubckt_1539_a3_x2 2 1116 1 1181 1186 88 a3_x2
xsubckt_1741_mx2_x2 1 1847 2 903 920 149 mx2_x2
xsubckt_1742_mx2_x2 1 1846 2 903 926 148 mx2_x2
xsubckt_118_mx2_x2 1 802 2 903 844 845 mx2_x2
xsubckt_653_oa22_x2 1 236 2 249 550 884 oa22_x2
xsubckt_663_o2_x2 1 227 2 256 863 o2_x2
xsubckt_821_nand3_x0 2 1 1709 1767 1775 45 nand3_x0
xsubckt_962_nand2_x0 2 1 1615 648 110 nand2_x0
xsubckt_995_nand4_x0 2 1 1590 620 742 747 761 nand4_x0
xsubckt_337_nand4_x0 2 1 544 680 691 708 793 nand4_x0
xsubckt_388_nand3_x0 2 1 493 784 833 20 nand3_x0
xsubckt_604_nand2_x0 2 1 284 566 661 nand2_x0
xsubckt_1299_nand3_x0 2 1 1343 773 780 164 nand3_x0
xsubckt_1343_a2_x2 1 1303 2 1304 1308 a2_x2
xsubckt_1569_a3_x2 2 1086 1 698 793 49 a3_x2
xsubckt_1858_sff1_x4 2 206 1 1875 174 sff1_x4
xsubckt_1819_sff1_x4 2 209 1 1905 85 sff1_x4
xsubckt_1770_sff1_x4 2 205 1 178 27 sff1_x4
xsubckt_1744_mx2_x2 1 1844 2 903 927 146 mx2_x2
xsubckt_1743_mx2_x2 1 1845 2 903 925 147 mx2_x2
xfeed_379 2 1 decap_w0
xfeed_378 2 1 decap_w0
xfeed_377 2 1 decap_w0
xfeed_376 2 1 decap_w0
xfeed_375 2 1 decap_w0
xfeed_374 2 1 decap_w0
xfeed_373 2 1 decap_w0
xfeed_372 2 1 tie
xfeed_371 2 1 decap_w0
xfeed_370 2 1 decap_w0
xsubckt_727_nand4_x0 2 1 1794 1795 1796 1797 1798 nand4_x0
xsubckt_1330_oa22_x2 1 1315 2 146 1384 1316 oa22_x2
xsubckt_1358_mx2_x2 1 1860 2 904 1290 44 mx2_x2
xsubckt_1449_o4_x2 1 1205 2 1207 1208 1421 281 o4_x2
xsubckt_1637_a2_x2 1 1018 2 1020 1160 a2_x2
xsubckt_1667_a2_x2 1 988 2 989 993 a2_x2
xsubckt_1748_mx2_x2 1 1842 2 903 1193 157 mx2_x2
xsubckt_914_nxr2_x1 1631 2 1 1641 888 nxr2_x1
xsubckt_1326_nxr2_x1 1318 2 1 1320 1327 nxr2_x1
xsubckt_1766_sff1_x4 2 205 1 182 31 sff1_x4
xfeed_385 2 1 decap_w0
xfeed_384 2 1 decap_w0
xfeed_383 2 1 decap_w0
xfeed_382 2 1 decap_w0
xfeed_381 2 1 decap_w0
xfeed_380 2 1 decap_w0
xsubckt_547_nand4_x0 2 1 337 480 681 17 832 nand4_x0
xsubckt_1672_nand3_x0 2 1 983 1181 1186 93 nand3_x0
xcmpt_abc_11873_new_n656_hfns_2 2 1 551 548 buf_x4
xcmpt_abc_11873_new_n656_hfns_1 2 1 548 549 buf_x4
xcmpt_abc_11873_new_n656_hfns_0 2 1 548 550 buf_x4
xsubckt_1545_nand2_x0 2 1 1110 1113 1160 nand2_x0
xsubckt_582_a4_x2 1 303 2 407 409 430 432 a4_x2
xsubckt_542_a4_x2 1 341 2 342 347 411 433 a4_x2
xsubckt_415_a3_x2 2 466 1 467 503 506 a3_x2
xsubckt_367_nand4_x0 2 1 514 691 708 831 27 nand4_x0
xsubckt_347_a4_x2 1 534 2 535 538 540 544 a4_x2
xsubckt_281_nand3_x0 2 1 603 681 697 713 nand3_x0
xsubckt_710_nand4_x0 2 1 1810 1812 1813 1814 1815 nand4_x0
xsubckt_988_nand3_x0 2 1 1596 461 612 761 nand3_x0
xsubckt_592_a4_x2 1 294 2 364 365 397 398 a4_x2
xsubckt_445_a3_x2 2 437 1 438 741 747 a3_x2
xsubckt_435_a3_x2 2 447 1 480 831 27 a3_x2
xsubckt_191_a3_x2 2 703 1 788 835 31 a3_x2
xsubckt_671_nand3_x0 2 1 220 262 269 134 nand3_x0
xsubckt_826_a4_x2 1 1704 2 1705 1706 1708 1785 a4_x2
xsubckt_553_a2_x2 1 331 2 332 333 a2_x2
xsubckt_358_a2_x2 1 523 2 524 529 a2_x2
xsubckt_729_a3_x2 2 1793 1 283 290 633 a3_x2
xsubckt_896_oa22_x2 1 1646 2 1655 1650 1651 oa22_x2
xsubckt_1134_nand3_x0 2 1 1481 1482 1484 1485 nand3_x0
xsubckt_1269_oa22_x2 1 1370 2 1380 579 877 oa22_x2
xsubckt_1275_nand2_x0 2 1 1364 1366 1370 nand2_x0
xsubckt_1665_nand2_x0 2 1 990 991 1160 nand2_x0
xsubckt_1575_nand2_x0 2 1 1080 1081 1087 nand2_x0
xsubckt_1302_ao22_x2 1 1340 2 891 1385 1342 ao22_x2
xsubckt_573_a2_x2 1 311 2 312 313 a2_x2
xsubckt_368_a2_x2 1 513 2 515 681 a2_x2
xsubckt_881_nand3_x0 2 1 1659 154 160 158 nand3_x0
xsubckt_971_nand3_x0 2 1 1608 1609 1614 620 nand3_x0
xsubckt_994_a3_x2 2 1591 1 742 746 761 a3_x2
xsubckt_1044_nand3_x0 2 1 1548 1549 1550 456 nand3_x0
xsubckt_1210_a4_x2 1 1412 2 1413 1414 1416 1427 a4_x2
xsubckt_1485_nand2_x0 2 1 1169 1171 1226 nand2_x0
xsubckt_397_nand4_x0 2 1 484 784 794 833 20 nand4_x0
xsubckt_184_nand2_x0 2 1 710 17 832 nand2_x0
xsubckt_242_oa22_x2 1 642 2 771 769 644 oa22_x2
xsubckt_1882_sff1_x4 2 202 1 1851 153 sff1_x4
xsubckt_1733_ao22_x2 1 1852 2 923 929 1151 ao22_x2
xsubckt_122_nor2_x0 2 1 796 17 27 nor2_x0
xsubckt_1046_a2_x2 1 1547 2 648 36 a2_x2
xsubckt_823_nand3_x0 2 1 1707 1773 577 700 nand3_x0
xsubckt_306_nand2_x0 2 1 578 580 680 nand2_x0
xsubckt_394_nand2_x0 2 1 487 488 489 nand2_x0
xsubckt_634_oa22_x2 1 254 2 486 568 878 oa22_x2
xsubckt_1622_a3_x2 2 1033 1 1181 1186 91 a3_x2
xsubckt_1843_sff1_x4 2 206 1 1889 66 sff1_x4
xsubckt_1804_sff1_x4 2 209 1 1920 61 sff1_x4
xsubckt_733_nand3_x0 2 1 1789 1791 559 583 nand3_x0
xsubckt_290_nand4_x0 2 1 594 691 832 23 834 nand4_x0
xsubckt_253_nand3_x0 2 1 631 680 698 718 nand3_x0
xsubckt_185_oa22_x2 1 709 2 710 715 723 oa22_x2
xsubckt_1403_oa22_x2 1 1248 2 1269 1260 1251 oa22_x2
xsubckt_1487_a3_x2 2 1167 1 591 793 113 a3_x2
xsubckt_1683_mx3_x2 2 1 972 1226 1146 1007 973 978 mx3_x2
xsubckt_1684_mx3_x2 2 1 971 1226 1146 1008 974 977 mx3_x2
xsubckt_1751_sff1_x4 2 208 1 1966 143 sff1_x4
xsubckt_1790_sff1_x4 2 210 1 1934 104 sff1_x4
xsubckt_1839_sff1_x4 2 211 1 1893 73 sff1_x4
xsubckt_1878_sff1_x4 2 207 1 1855 53 sff1_x4
xsubckt_1167_mx2_x2 1 1888 2 1460 11 1453 mx2_x2
xsubckt_1166_mx2_x2 1 1453 2 1458 1454 1455 mx2_x2
xsubckt_1165_mx2_x2 1 1454 2 585 92 152 mx2_x2
xsubckt_784_nand2_x0 2 1 1741 1742 1743 nand2_x0
xsubckt_1337_nand2_x0 2 1 1309 1379 45 nand2_x0
xsubckt_1464_nand3_x0 2 1 1190 1191 1773 671 nand3_x0
xsubckt_1477_oa22_x2 1 1177 2 1773 671 869 oa22_x2
xsubckt_1307_nxr2_x1 1335 2 1 1338 1345 nxr2_x1
xsubckt_1786_sff1_x4 2 206 1 1937 122 sff1_x4
xcmpt_abc_11873_new_n504_hfns_3 2 1 720 716 buf_x4
xcmpt_abc_11873_new_n504_hfns_2 2 1 716 717 buf_x4
xcmpt_abc_11873_new_n504_hfns_1 2 1 716 718 buf_x4
xcmpt_abc_11873_new_n504_hfns_0 2 1 716 719 buf_x4
xcmpt_abc_11873_new_n506_hfns_2 2 1 714 711 buf_x4
xcmpt_abc_11873_new_n506_hfns_1 2 1 711 712 buf_x4
xcmpt_abc_11873_new_n506_hfns_0 2 1 711 713 buf_x4
xsubckt_1067_nand2_x0 2 1 1533 647 829 nand2_x0
xsubckt_1016_nand3_x0 2 1 1569 1572 1593 1596 nand3_x0
xsubckt_776_ao22_x2 1 1748 2 1776 1784 151 ao22_x2
xsubckt_215_a4_x2 1 672 2 787 792 25 836 a4_x2
xsubckt_156_nand2_x0 2 1 748 750 751 nand2_x0
xsubckt_539_a4_x2 1 344 2 345 346 518 520 a4_x2
xsubckt_1293_oa22_x2 1 1348 2 150 1384 1349 oa22_x2
xsubckt_1457_nand2_x0 2 1 1197 1199 1233 nand2_x0
xsubckt_1215_oa22_x2 1 1407 2 715 710 569 oa22_x2
xsubckt_0_inv_x0 2 1 83 917 inv_x0
xsubckt_1_inv_x0 2 1 71 916 inv_x0
xsubckt_2_inv_x0 2 1 41 915 inv_x0
xsubckt_3_inv_x0 2 1 102 914 inv_x0
xsubckt_4_inv_x0 2 1 64 913 inv_x0
xsubckt_1050_nand2_x0 2 1 1545 648 82 nand2_x0
xsubckt_862_a3_x2 2 1674 1 1675 1676 1677 a3_x2
xsubckt_832_a3_x2 2 1699 1 1700 1701 1702 a3_x2
xsubckt_761_nor2_x0 2 1 1761 1762 1765 nor2_x0
xsubckt_315_nand3_x0 2 1 569 691 833 20 nand3_x0
xsubckt_256_a2_x2 1 628 2 629 774 a2_x2
xsubckt_189_nand4_x0 2 1 705 708 17 26 836 nand4_x0
xsubckt_5_inv_x0 2 1 36 912 inv_x0
xsubckt_6_inv_x0 2 1 12 911 inv_x0
xsubckt_7_inv_x0 2 1 110 910 inv_x0
xsubckt_8_inv_x0 2 1 42 909 inv_x0
xsubckt_9_inv_x0 2 1 39 908 inv_x0
xsubckt_405_nand3_x0 2 1 476 681 707 713 nand3_x0
xsubckt_431_a2_x2 1 451 2 452 457 a2_x2
xsubckt_493_nand3_x0 2 1 390 575 591 795 nand3_x0
xsubckt_950_a2_x2 1 1621 2 847 10 a2_x2
xsubckt_883_nand3_x0 2 1 1657 894 895 158 nand3_x0
xsubckt_882_a3_x2 2 1658 1 894 895 158 a3_x2
xsubckt_750_oa22_x2 1 1772 2 719 688 515 oa22_x2
xsubckt_745_a2_x2 1 1777 2 1778 577 a2_x2
xsubckt_705_nand3_x0 2 1 1815 262 268 115 nand3_x0
xsubckt_286_nor3_x0 2 1 598 601 604 634 nor3_x0
xsubckt_491_a2_x2 1 391 2 392 508 a2_x2
xsubckt_1322_ao22_x2 1 1322 2 888 1385 1324 ao22_x2
xsubckt_901_mx2_x2 1 1642 2 562 89 149 mx2_x2
xsubckt_900_mx2_x2 1 1965 2 1662 142 1643 mx2_x2
xsubckt_742_nand4_x0 2 1 1780 1783 593 664 686 nand4_x0
xsubckt_399_nand4_x0 2 1 482 483 485 488 489 nand4_x0
xsubckt_1499_nor4_x0 2 1 1155 1160 1167 1168 289 nor4_x0
xsubckt_1593_oa22_x2 1 1062 2 218 1205 1064 oa22_x2
xsubckt_1219_nand2_x0 2 1 1403 1404 539 nand2_x0
xsubckt_1041_a3_x2 2 1551 1 456 741 749 a3_x2
xsubckt_902_mx2_x2 1 1964 2 1662 141 1642 mx2_x2
xsubckt_254_mx3_x2 2 1 630 916 9 840 841 842 mx3_x2
xsubckt_1397_nand2_x0 2 1 1254 580 148 nand2_x0
xsubckt_1554_oa22_x2 1 1101 2 1820 1205 1103 oa22_x2
xsubckt_1714_ao22_x2 1 941 2 950 943 942 ao22_x2
xsubckt_1824_sff1_x4 2 211 1 91 99 sff1_x4
xsubckt_1863_sff1_x4 2 206 1 1870 169 sff1_x4
xsubckt_1535_mx3_x2 2 1 1120 1226 1129 1194 1126 1123 mx3_x2
xsubckt_1534_mx3_x2 2 1 1121 1226 1128 1193 1122 1127 mx3_x2
xsubckt_1405_mx2_x2 1 1856 2 903 1247 54 mx2_x2
xsubckt_699_nand4_x0 2 1 1820 1823 1824 1825 1826 nand4_x0
xsubckt_966_nand2_x0 2 1 1612 648 39 nand2_x0
xsubckt_1080_nand2_x0 2 1 1521 1543 1587 nand2_x0
xsubckt_1142_mx3_x2 2 1 1474 585 445 807 108 893 mx3_x2
xsubckt_1208_a2_x2 1 1414 2 1415 706 a2_x2
xsubckt_1859_sff1_x4 2 206 1 1874 173 sff1_x4
xsubckt_1697_nand2_x0 2 1 958 990 992 nand2_x0
xsubckt_1669_a3_x2 2 986 1 698 793 59 a3_x2
xsubckt_1649_a3_x2 2 1006 1 698 793 58 a3_x2
xsubckt_1463_a2_x2 1 1191 2 663 777 a2_x2
xsubckt_1462_oa22_x2 1 1192 2 1773 671 870 oa22_x2
xsubckt_1423_a2_x2 1 1230 2 1231 1236 a2_x2
xsubckt_382_nand4_x0 2 1 499 610 612 645 767 nand4_x0
xsubckt_131_oa22_x2 1 773 2 917 177 64 oa22_x2
xsubckt_814_ao22_x2 1 1715 2 1776 1784 146 ao22_x2
xsubckt_1076_nand3_x0 2 1 1524 1525 1528 1583 nand3_x0
xsubckt_1225_o4_x2 1 1397 2 1398 1417 1782 554 o4_x2
xsubckt_1265_ao22_x2 1 1373 2 1374 1376 1388 ao22_x2
xsubckt_1771_sff1_x4 2 210 1 1952 137 sff1_x4
xsubckt_1727_a2_x2 1 928 2 1144 1156 a2_x2
xsubckt_1717_a2_x2 1 938 2 939 1069 a2_x2
xsubckt_1288_a2_x2 1 1352 2 1353 1354 a2_x2
xsubckt_645_nand3_x0 2 1 244 262 269 136 nand3_x0
xsubckt_689_oa22_x2 1 1829 2 486 568 874 oa22_x2
xsubckt_786_nand2_x0 2 1 1739 1740 1745 nand2_x0
xsubckt_1173_ao22_x2 1 1447 2 1449 1452 585 ao22_x2
xsubckt_1202_nand2_x0 2 1 1420 1438 475 nand2_x0
xsubckt_1767_sff1_x4 2 205 1 181 30 sff1_x4
xsubckt_1680_nand2_x0 2 1 975 976 977 nand2_x0
xsubckt_1618_ao22_x2 1 1037 2 230 1206 1039 ao22_x2
xsubckt_1331_oa22_x2 1 1314 2 46 1377 1315 oa22_x2
xsubckt_1286_nand3_x0 2 1 1354 1356 1364 1373 nand3_x0
xsubckt_10_inv_x0 2 1 159 907 inv_x0
xsubckt_11_inv_x0 2 1 106 906 inv_x0
xsubckt_12_inv_x0 2 1 9 905 inv_x0
xsubckt_13_inv_x0 2 1 4 900 inv_x0
xsubckt_14_inv_x0 2 1 107 899 inv_x0
xsubckt_1022_nand2_x0 2 1 1564 1565 1567 nand2_x0
xsubckt_375_nand3_x0 2 1 506 681 707 719 nand3_x0
xsubckt_15_inv_x0 2 1 109 898 inv_x0
xsubckt_16_inv_x0 2 1 153 897 inv_x0
xsubckt_17_inv_x0 2 1 152 896 inv_x0
xsubckt_18_inv_x0 2 1 160 895 inv_x0
xsubckt_19_inv_x0 2 1 154 894 inv_x0
xsubckt_163_a4_x2 1 738 2 741 749 755 760 a4_x2
xsubckt_234_ao22_x2 1 653 2 654 660 800 ao22_x2
xsubckt_757_ao22_x2 1 1765 2 1776 1784 153 ao22_x2
xsubckt_796_ao22_x2 1 1731 2 1827 1822 1792 ao22_x2
xsubckt_915_nxr2_x1 1630 2 1 1631 1636 nxr2_x1
xsubckt_996_nand2_x0 2 1 1589 1590 739 nand2_x0
xsubckt_1069_nand2_x0 2 1 1531 1532 1575 nand2_x0
xsubckt_1586_nand3_x0 2 1 1069 1070 1075 1090 nand3_x0
xsubckt_1526_ao22_x2 1 1129 2 1811 1206 1131 ao22_x2
xsubckt_501_nand2_x0 2 1 382 730 766 nand2_x0
xsubckt_466_nxr2_x1 416 2 1 417 885 nxr2_x1
xsubckt_765_nand3_x0 2 1 1758 1767 1775 58 nand3_x0
xsubckt_1496_nand3_x0 2 1 1158 1160 1162 1163 nand3_x0
xsubckt_142_ao22_x2 1 762 2 71 91 774 ao22_x2
xsubckt_134_a2_x2 1 770 2 771 774 a2_x2
xsubckt_124_a2_x2 1 789 2 22 20 a2_x2
xsubckt_269_ao22_x2 1 615 2 622 626 628 ao22_x2
xsubckt_284_nor4_x0 2 1 600 601 636 641 651 nor4_x0
xsubckt_672_a4_x2 1 219 2 220 221 222 223 a4_x2
xsubckt_897_nxr2_x1 1645 2 1 1658 150 nxr2_x1
xsubckt_555_a3_x2 2 329 1 330 345 346 a3_x2
xsubckt_317_nand3_x0 2 1 567 570 681 713 nand3_x0
xsubckt_770_a3_x2 2 1753 1 1754 1757 1758 a3_x2
xsubckt_801_nand2_x0 2 1 1726 1727 1728 nand2_x0
xsubckt_1666_oa22_x2 1 989 2 1160 991 1155 oa22_x2
xsubckt_1627_oa22_x2 1 1028 2 1032 1034 1188 oa22_x2
xsubckt_488_a2_x2 1 394 2 395 400 a2_x2
xsubckt_354_nand4_x0 2 1 527 787 832 835 31 nand4_x0
xsubckt_707_nand3_x0 2 1 1813 262 269 131 nand3_x0
xsubckt_731_oa22_x2 1 1791 2 496 565 790 oa22_x2
xsubckt_777_nor2_x0 2 1 1747 1748 1749 nor2_x0
xsubckt_848_nand2_x0 2 1 1686 1780 89 nand2_x0
xsubckt_907_a2_x2 1 1637 2 1638 1640 a2_x2
xsubckt_1182_oa22_x2 1 1440 2 494 713 780 oa22_x2
xsubckt_1380_a4_x2 1 1269 2 1270 1282 1291 1300 a4_x2
xsubckt_1377_ao22_x2 1 1272 2 806 1387 1273 ao22_x2
xsubckt_563_o3_x2 1 321 2 492 677 832 o3_x2
xsubckt_351_nand2_x0 2 1 530 658 793 nand2_x0
xsubckt_300_nand3_x0 2 1 584 597 680 718 nand3_x0
xsubckt_654_nand4_x0 2 1 235 236 237 238 239 nand4_x0
xsubckt_997_a2_x2 1 1588 2 1589 1609 a2_x2
xsubckt_1883_sff1_x4 2 202 1 1850 152 sff1_x4
xsubckt_1844_sff1_x4 2 209 1 1888 11 sff1_x4
xsubckt_1805_sff1_x4 2 205 1 1919 60 sff1_x4
xsubckt_1602_mx2_x2 1 1053 2 1227 1054 1087 mx2_x2
xsubckt_1601_mx2_x2 1 1054 2 1063 1055 1057 mx2_x2
xsubckt_1537_a3_x2 2 1118 1 698 793 48 a3_x2
xsubckt_1511_nand3_x0 2 1 1144 1153 1169 1210 nand3_x0
xsubckt_486_o2_x2 1 396 2 541 677 o2_x2
xsubckt_477_ao22_x2 1 405 2 761 740 755 ao22_x2
xsubckt_831_nand2_x0 2 1 1700 1769 152 nand2_x0
xsubckt_968_nand2_x0 2 1 1929 1611 1612 nand2_x0
xsubckt_1068_a3_x2 2 1532 1 755 760 767 a3_x2
xsubckt_1082_nand2_x0 2 1 1519 1578 650 nand2_x0
xsubckt_1211_ao22_x2 1 1411 2 1429 1419 1412 ao22_x2
xsubckt_1263_a3_x2 2 1375 1 773 780 168 a3_x2
xsubckt_1879_sff1_x4 2 207 1 1854 52 sff1_x4
xsubckt_1642_ao22_x2 1 1013 2 1203 1789 152 ao22_x2
xsubckt_1605_a2_x2 1 1050 2 1052 1160 a2_x2
xsubckt_350_ao22_x2 1 531 2 642 532 533 ao22_x2
xsubckt_294_nand4_x0 2 1 590 22 834 835 31 nand4_x0
xsubckt_674_oa22_x2 1 217 2 486 568 875 oa22_x2
xsubckt_1047_oa22_x2 1 1914 2 1559 1558 1547 oa22_x2
xsubckt_1207_ao22_x2 1 1415 2 17 590 527 ao22_x2
xsubckt_1791_sff1_x4 2 211 1 1933 103 sff1_x4
xsubckt_1752_sff1_x4 2 207 1 1965 142 sff1_x4
xsubckt_1292_nand2_x0 2 1 1349 1350 550 nand2_x0
xsubckt_414_nor4_x0 2 1 467 468 472 482 490 nor4_x0
xsubckt_647_nand3_x0 2 1 242 263 268 128 nand3_x0
xsubckt_788_nand2_x0 2 1 1738 1792 1833 nand2_x0
xsubckt_1176_mx2_x2 1 1444 2 586 1445 93 mx2_x2
xsubckt_1222_nor4_x0 2 1 1400 1401 1402 1405 1408 nor4_x0
xsubckt_1787_sff1_x4 2 209 1 1936 64 sff1_x4
xsubckt_1685_a2_x2 1 970 2 972 979 a2_x2
xsubckt_1677_ao22_x2 1 978 2 984 986 1189 ao22_x2
xsubckt_1347_nxr2_x1 1299 2 1 1302 1313 nxr2_x1
xsubckt_781_ao22_x2 1 1744 2 1776 1784 150 ao22_x2
xsubckt_1024_nand2_x0 2 1 1563 647 868 nand2_x0
xsubckt_1061_nand3_x0 2 1 1537 1538 1585 1619 nand3_x0
xsubckt_1154_ao22_x2 1 1464 2 1465 1466 1467 ao22_x2
xsubckt_1177_mx2_x2 1 1887 2 1446 1444 111 mx2_x2
xsubckt_1178_mx2_x2 1 1886 2 9 113 192 mx2_x2
xsubckt_1704_nxr2_x1 951 2 1 952 1044 nxr2_x1
xsubckt_1451_nand3_x0 2 1 1203 530 568 585 nand3_x0
xsubckt_467_nand3_x0 2 1 415 698 719 800 nand3_x0
xsubckt_377_nand3_x0 2 1 504 612 617 753 nand3_x0
xsubckt_291_nand2_x0 2 1 593 595 17 nand2_x0
xsubckt_720_nand3_x0 2 1 1801 262 268 114 nand3_x0
xsubckt_771_nand2_x0 2 1 1983 1753 1759 nand2_x0
xsubckt_861_nand2_x0 2 1 1675 1769 147 nand2_x0
xcmpt_abc_11873_new_n518_hfns_2 2 1 699 696 buf_x4
xcmpt_abc_11873_new_n518_hfns_1 2 1 696 697 buf_x4
xcmpt_abc_11873_new_n518_hfns_0 2 1 696 698 buf_x4
xsubckt_1643_o2_x2 1 1012 2 1200 808 o2_x2
xsubckt_1546_ao22_x2 1 1109 2 1161 1112 1154 ao22_x2
xsubckt_1488_o2_x2 1 1166 2 1168 289 o2_x2
xsubckt_1361_nand3_x0 2 1 1287 773 780 174 nand3_x0
xsubckt_630_nand3_x0 2 1 258 263 269 145 nand3_x0
xsubckt_503_nand2_x0 2 1 380 382 460 nand2_x0
xsubckt_355_a4_x2 1 526 2 788 794 835 31 a4_x2
xsubckt_335_a4_x2 1 546 2 547 552 556 558 a4_x2
xsubckt_1023_ao22_x2 1 1921 2 1574 1564 1568 ao22_x2
xcmpt_abc_11873_new_n479_hfns_2 2 1 748 745 buf_x4
xcmpt_abc_11873_new_n479_hfns_1 2 1 745 746 buf_x4
xcmpt_abc_11873_new_n479_hfns_0 2 1 745 747 buf_x4
xsubckt_1493_ao22_x2 1 1161 2 1772 672 60 ao22_x2
xsubckt_590_a4_x2 1 296 2 491 495 582 584 a4_x2
xsubckt_450_nand3_x0 2 1 432 528 680 17 nand3_x0
xsubckt_413_nand2_x0 2 1 468 469 470 nand2_x0
xsubckt_1144_nand2_x0 2 1 1891 1473 1475 nand2_x0
xsubckt_1271_nand3_x0 2 1 1368 566 794 915 nand3_x0
xsubckt_1216_oa22_x2 1 1406 2 715 710 695 oa22_x2
xsubckt_981_nand2_x0 2 1 1925 1602 1603 nand2_x0
xsubckt_932_a3_x2 2 1623 1 1663 262 269 a3_x2
xsubckt_1583_nor3_x0 2 1 1072 1073 1074 1161 nor3_x0
xsubckt_1454_ao22_x2 1 1200 2 790 695 514 ao22_x2
xsubckt_531_a2_x2 1 352 2 353 354 a2_x2
xsubckt_360_nand3_x0 2 1 521 658 17 832 nand3_x0
xsubckt_336_a2_x2 1 545 2 546 560 a2_x2
xsubckt_737_a3_x2 2 1785 1 1786 1788 1790 a3_x2
xsubckt_840_nand3_x0 2 1 1693 1767 1775 56 nand3_x0
xsubckt_891_nand2_x0 2 1 1650 1659 893 nand2_x0
xsubckt_1003_a4_x2 1 1582 2 1585 1587 627 753 a4_x2
xsubckt_977_nand3_x0 2 1 1604 1614 614 620 nand3_x0
xsubckt_797_a3_x2 2 1730 1 1767 1775 48 a3_x2
xsubckt_100_inv_x0 2 1 77 813 inv_x0
xsubckt_101_inv_x0 2 1 97 812 inv_x0
xsubckt_102_inv_x0 2 1 195 811 inv_x0
xsubckt_103_inv_x0 2 1 76 810 inv_x0
xsubckt_105_inv_x0 2 1 809 93 inv_x0
xsubckt_158_ao22_x2 1 743 2 71 92 774 ao22_x2
xsubckt_356_nand4_x0 2 1 525 788 793 835 31 nand4_x0
xsubckt_1073_a4_x2 1 1527 2 1541 378 753 767 a4_x2
xsubckt_712_oa22_x2 1 1808 2 253 700 888 oa22_x2
xsubckt_246_o3_x2 1 638 2 639 683 686 o3_x2
xsubckt_107_inv_x0 2 1 808 92 inv_x0
xsubckt_109_inv_x0 2 1 807 91 inv_x0
xsubckt_1608_oa22_x2 1 1047 2 1160 1052 1155 oa22_x2
xsubckt_1250_nand4_x0 2 1 1388 1389 1391 1783 390 nand4_x0
xsubckt_1101_a3_x2 2 1504 1 1515 1541 746 a3_x2
xsubckt_1083_a4_x2 1 1518 2 1521 1522 1578 650 a4_x2
xsubckt_911_mx2_x2 1 1963 2 1662 140 1634 mx2_x2
xsubckt_910_mx2_x2 1 1634 2 563 1635 88 mx2_x2
xsubckt_302_nand3_x0 2 1 582 591 718 799 nand3_x0
xsubckt_139_o2_x2 1 765 2 91 70 o2_x2
xsubckt_480_nand3_x0 2 1 402 497 792 800 nand3_x0
xsubckt_1171_a3_x2 2 1449 1 1450 1451 908 a3_x2
xsubckt_1004_a2_x2 1 1581 2 1609 766 a2_x2
xsubckt_917_mx2_x2 1 1962 2 1662 139 1629 mx2_x2
xsubckt_916_mx2_x2 1 1629 2 563 1630 87 mx2_x2
xsubckt_833_nand2_x0 2 1 1969 1699 1703 nand2_x0
xsubckt_803_o2_x2 1 1724 2 1725 1730 o2_x2
xsubckt_1387_a4_x2 1 1263 2 1264 1265 1266 550 a4_x2
xsubckt_1424_nxr2_x1 1229 2 1 1230 1238 nxr2_x1
xsubckt_1513_nand3_x0 2 1 1142 697 795 47 nand3_x0
xsubckt_1620_a3_x2 2 1035 1 697 795 51 a3_x2
xsubckt_1654_nand2_x0 2 1 1001 1003 1005 nand2_x0
xsubckt_1715_ao22_x2 1 940 2 1091 1076 1071 ao22_x2
xsubckt_1825_sff1_x4 2 211 1 90 98 sff1_x4
xsubckt_1864_sff1_x4 2 202 1 1869 59 sff1_x4
xsubckt_1029_nand4_x0 2 1 1560 1561 378 609 621 nand4_x0
xsubckt_1026_mx2_x2 1 1919 2 648 1567 60 mx2_x2
xsubckt_780_nand3_x0 2 1 1745 1767 1775 50 nand3_x0
xsubckt_655_oa22_x2 1 190 2 288 240 235 oa22_x2
xsubckt_370_ao22_x2 1 511 2 911 652 512 ao22_x2
xsubckt_1333_nand3_x0 2 1 1312 1314 1319 1327 nand3_x0
xsubckt_1416_mx2_x2 1 1855 2 904 1237 53 mx2_x2
xsubckt_1495_a3_x2 2 1159 1 1160 1162 1163 a3_x2
xsubckt_1500_o4_x2 1 1154 2 1160 1167 1168 289 o4_x2
xsubckt_1203_nor4_x0 2 1 1419 1420 1421 1439 1787 nor4_x0
xsubckt_879_mx2_x2 1 1968 2 1662 145 1661 mx2_x2
xsubckt_878_mx2_x2 1 1661 2 562 93 153 mx2_x2
xsubckt_512_nand3_x0 2 1 371 612 618 753 nand3_x0
xsubckt_1371_mx2_x2 1 1859 2 904 1278 57 mx2_x2
xsubckt_1378_a2_x2 1 1271 2 1272 1277 a2_x2
xsubckt_1498_oa22_x2 1 1156 2 1210 1169 1159 oa22_x2
xsubckt_1772_sff1_x4 2 208 1 1951 136 sff1_x4
xsubckt_920_nxr2_x1 1626 2 1 1627 1628 nxr2_x1
xsubckt_20_inv_x0 2 1 151 893 inv_x0
xsubckt_21_inv_x0 2 1 150 892 inv_x0
xsubckt_596_nand4_x0 2 1 178 291 300 301 352 nand4_x0
xsubckt_1459_oa22_x2 1 1195 2 146 1201 1197 oa22_x2
xsubckt_863_nand2_x0 2 1 1978 1674 1678 nand2_x0
xsubckt_22_inv_x0 2 1 149 891 inv_x0
xsubckt_23_inv_x0 2 1 148 890 inv_x0
xsubckt_24_inv_x0 2 1 155 889 inv_x0
xsubckt_25_inv_x0 2 1 147 888 inv_x0
xsubckt_26_inv_x0 2 1 146 887 inv_x0
xsubckt_559_oa22_x2 1 325 2 375 379 644 oa22_x2
xsubckt_1768_sff1_x4 2 205 1 180 29 sff1_x4
xsubckt_1043_ao22_x2 1 1549 2 732 736 102 ao22_x2
xsubckt_293_a4_x2 1 591 2 23 834 835 31 a4_x2
xsubckt_238_nand4_x0 2 1 649 783 788 793 9 nand4_x0
xsubckt_27_inv_x0 2 1 108 886 inv_x0
xsubckt_28_inv_x0 2 1 105 885 inv_x0
xsubckt_29_inv_x0 2 1 11 884 inv_x0
xsubckt_126_a3_x2 2 781 1 783 787 794 a3_x2
xsubckt_1566_ao22_x2 1 1089 2 805 1200 1265 ao22_x2
xsubckt_567_a4_x2 1 317 2 318 325 326 347 a4_x2
xsubckt_577_a4_x2 1 308 2 535 538 666 669 a4_x2
xsubckt_587_a4_x2 1 299 2 425 426 477 481 a4_x2
xsubckt_898_nxr2_x1 1644 2 1 1645 1646 nxr2_x1
xsubckt_850_a3_x2 2 1684 1 1685 1686 1687 a3_x2
xsubckt_805_nand2_x0 2 1 1723 1792 1810 nand2_x0
xsubckt_214_a2_x2 1 673 2 674 676 a2_x2
xsubckt_325_nand2_x0 2 1 559 570 718 nand2_x0
xsubckt_1536_nand2_x0 2 1 1119 1121 1134 nand2_x0
xsubckt_880_a3_x2 2 1660 1 154 160 158 a3_x2
xsubckt_743_nor2_x0 2 1 1779 474 660 nor2_x0
xsubckt_274_a2_x2 1 610 2 754 760 a2_x2
xsubckt_1446_nand2_x0 2 1 1208 1438 539 nand2_x0
xsubckt_1089_nand4_x0 2 1 1513 1575 378 753 767 nand4_x0
xsubckt_793_a2_x2 1 1733 2 1734 1735 a2_x2
xsubckt_418_o3_x2 1 183 2 464 599 604 o3_x2
xsubckt_588_a2_x2 1 298 2 299 319 a2_x2
xsubckt_1304_ao22_x2 1 1338 2 874 1378 1340 ao22_x2
xsubckt_1356_nand2_x0 2 1 1291 1293 1298 nand2_x0
xsubckt_1410_a4_x2 1 1242 2 1243 1244 1245 550 a4_x2
xsubckt_1125_nand3_x0 2 1 1490 1668 899 907 nand3_x0
xsubckt_767_oa22_x2 1 1756 2 1770 1771 855 oa22_x2
xsubckt_728_oa22_x2 1 184 2 288 1799 1794 oa22_x2
xsubckt_1810_sff1_x4 2 211 1 1914 36 sff1_x4
xsubckt_1212_ao22_x2 1 1410 2 570 698 719 ao22_x2
xsubckt_1098_nor2_x0 2 1 1904 1506 1510 nor2_x0
xsubckt_1086_nand2_x0 2 1 1516 647 828 nand2_x0
xsubckt_1035_nand3_x0 2 1 1556 615 730 740 nand3_x0
xsubckt_835_nand2_x0 2 1 1697 1707 174 nand2_x0
xsubckt_711_o2_x2 1 1809 2 256 858 o2_x2
xsubckt_392_nand3_x0 2 1 489 497 681 713 nand3_x0
xsubckt_533_nor3_x0 2 1 350 14 155 12 nor3_x0
xsubckt_1290_ao22_x2 1 1351 2 1379 580 50 ao22_x2
xsubckt_1515_nand3_x0 2 1 1140 1181 1186 87 nand3_x0
xsubckt_1611_mx2_x2 1 1044 2 1053 1048 1050 mx2_x2
xsubckt_1612_mx2_x2 1 1043 2 1053 1047 1049 mx2_x2
xsubckt_1693_nand3_x0 2 1 962 963 966 969 nand3_x0
xsubckt_1884_sff1_x4 2 202 1 1849 151 sff1_x4
xsubckt_1256_a2_x2 1 1382 2 1383 777 a2_x2
xsubckt_1247_ao22_x2 1 1391 2 777 773 721 ao22_x2
xsubckt_1206_a2_x2 1 1416 2 1418 1783 a2_x2
xsubckt_439_ao22_x2 1 443 2 543 688 719 ao22_x2
xsubckt_636_oa22_x2 1 252 2 542 702 715 oa22_x2
xsubckt_1806_sff1_x4 2 209 1 1918 40 sff1_x4
xsubckt_1845_sff1_x4 2 208 1 1887 111 sff1_x4
xsubckt_1229_mx2_x2 1 1885 2 1394 1984 168 mx2_x2
xsubckt_551_nand4_x0 2 1 333 480 681 831 27 nand4_x0
xsubckt_1386_nand2_x0 2 1 1264 580 149 nand2_x0
xsubckt_1391_nxr2_x1 1259 2 1 1261 1269 nxr2_x1
xsubckt_1735_a2_x2 1 921 2 922 962 a2_x2
xsubckt_1753_sff1_x4 2 207 1 1964 141 sff1_x4
xsubckt_1792_sff1_x4 2 210 1 1932 42 sff1_x4
xsubckt_1014_nand4_x0 2 1 1571 627 729 742 747 nand4_x0
xsubckt_955_nand2_x0 2 1 1620 647 42 nand2_x0
xsubckt_904_nand3_x0 2 1 1640 155 160 158 nand3_x0
xsubckt_334_nand3_x0 2 1 547 566 794 799 nand3_x0
xsubckt_598_nand4_x0 2 1 289 290 486 564 568 nand4_x0
xsubckt_1576_mx2_x2 1 1079 2 1082 1176 1189 mx2_x2
xsubckt_1065_nand3_x0 2 1 1534 1535 408 737 nand3_x0
xsubckt_865_nand2_x0 2 1 1672 1707 169 nand2_x0
xsubckt_775_nand2_x0 2 1 1749 1750 1751 nand2_x0
xsubckt_295_nand2_x0 2 1 589 591 713 nand2_x0
xsubckt_1313_oa22_x2 1 1330 2 148 1384 1332 oa22_x2
xsubckt_1551_ao22_x2 1 1104 2 890 1202 1106 ao22_x2
xsubckt_1590_ao22_x2 1 1065 2 892 1202 1067 ao22_x2
xsubckt_1639_ao22_x2 1 1016 2 1161 1019 1154 ao22_x2
xsubckt_1686_nand2_x0 2 1 969 972 979 nand2_x0
xsubckt_1749_sff1_x4 2 208 1 1968 145 sff1_x4
xsubckt_1788_sff1_x4 2 205 1 10 65 sff1_x4
xsubckt_1508_o2_x2 1 1147 2 1148 1150 o2_x2
xsubckt_1548_o2_x2 1 1107 2 1200 804 o2_x2
xsubckt_1705_nxr2_x1 950 2 1 952 1043 nxr2_x1
xsubckt_1267_nor2_x0 2 1 1371 1372 1373 nor2_x0
xsubckt_709_a4_x2 1 1811 2 1812 1813 1814 1815 a4_x2
xsubckt_660_a4_x2 1 230 2 231 232 233 234 a4_x2
xsubckt_338_a3_x2 2 543 1 708 835 31 a3_x2
xsubckt_513_a3_x2 2 370 1 371 372 373 a3_x2
xsubckt_544_nand3_x0 2 1 181 340 356 367 nand3_x0
xsubckt_1007_nand3_x0 2 1 1578 1580 378 753 nand3_x0
xsubckt_807_nand2_x0 2 1 1721 1774 147 nand2_x0
xsubckt_223_nand4_x0 2 1 664 708 832 26 836 nand4_x0
xsubckt_132_a2_x2 1 772 2 810 71 a2_x2
xsubckt_543_a3_x2 2 340 1 341 600 605 a3_x2
xsubckt_583_a3_x2 2 302 1 303 304 334 a3_x2
xsubckt_608_ao22_x2 1 280 2 831 527 492 ao22_x2
xsubckt_1095_nand3_x0 2 1 1508 1543 1587 753 nand3_x0
xsubckt_877_a3_x2 2 1662 1 1663 263 269 a3_x2
xsubckt_703_nand4_x0 2 1 1816 1817 1818 1819 248 nand4_x0
xsubckt_111_inv_x0 2 1 806 90 inv_x0
xsubckt_400_nand2_x0 2 1 481 660 680 nand2_x0
xsubckt_476_a2_x2 1 406 2 407 409 a2_x2
xsubckt_613_nand4_x0 2 1 275 276 282 777 33 nand4_x0
xsubckt_1311_nand2_x0 2 1 1332 1334 550 nand2_x0
xsubckt_1131_nand2_x0 2 1 1484 777 87 nand2_x0
xsubckt_791_oa22_x2 1 1735 2 1770 1771 852 oa22_x2
xsubckt_713_oa22_x2 1 1807 2 486 568 872 oa22_x2
xsubckt_249_nor3_x0 2 1 635 636 641 651 nor3_x0
xsubckt_113_inv_x0 2 1 805 89 inv_x0
xsubckt_115_inv_x0 2 1 804 88 inv_x0
xsubckt_117_inv_x0 2 1 803 87 inv_x0
xsubckt_496_a2_x2 1 387 2 388 504 a2_x2
xsubckt_574_nand3_x0 2 1 310 311 314 635 nand3_x0
xsubckt_1324_ao22_x2 1 1320 2 872 1378 1322 ao22_x2
xsubckt_1395_nand3_x0 2 1 1256 773 780 171 nand3_x0
xsubckt_1560_oa22_x2 1 1095 2 1098 1099 1175 oa22_x2
xsubckt_1648_oa22_x2 1 1007 2 240 1205 1009 oa22_x2
xsubckt_1254_nand4_x0 2 1 1384 1783 577 593 709 nand4_x0
xsubckt_921_mx2_x2 1 1625 2 563 1626 86 mx2_x2
xsubckt_787_oa22_x2 1 1975 2 218 1792 1739 oa22_x2
xsubckt_119_inv_x0 2 1 802 86 inv_x0
xsubckt_447_nand2_x0 2 1 435 437 613 nand2_x0
xsubckt_484_nand3_x0 2 1 398 707 719 800 nand3_x0
xsubckt_1521_nand2_x0 2 1 1134 1136 1154 nand2_x0
xsubckt_1830_sff1_x4 2 210 1 1902 67 sff1_x4
xsubckt_1251_a3_x2 2 1387 1 1783 593 709 a3_x2
xsubckt_1074_nand4_x0 2 1 1526 1541 378 753 767 nand4_x0
xsubckt_1072_oa22_x2 1 1528 2 1529 1531 611 oa22_x2
xsubckt_964_nand3_x0 2 1 1613 1614 355 620 nand3_x0
xsubckt_927_mx2_x2 1 1957 2 1624 118 1643 mx2_x2
xsubckt_926_mx2_x2 1 1958 2 1624 119 1647 mx2_x2
xsubckt_925_mx2_x2 1 1959 2 1624 120 1652 mx2_x2
xsubckt_924_mx2_x2 1 1960 2 1624 121 1661 mx2_x2
xsubckt_922_mx2_x2 1 1961 2 1662 138 1625 mx2_x2
xsubckt_837_nand2_x0 2 1 1695 1780 91 nand2_x0
xsubckt_259_o2_x2 1 625 2 88 71 o2_x2
xsubckt_424_ao22_x2 1 458 2 644 459 463 ao22_x2
xsubckt_610_nand2_x0 2 1 278 521 553 nand2_x0
xsubckt_1341_nand2_x0 2 1 1305 580 153 nand2_x0
xsubckt_1517_oa22_x2 1 1138 2 1140 1142 1165 oa22_x2
xsubckt_1556_oa22_x2 1 1099 2 1115 1117 1188 oa22_x2
xsubckt_1174_a2_x2 1 1446 2 1447 1448 a2_x2
xsubckt_1164_a2_x2 1 1455 2 1456 1457 a2_x2
xsubckt_1033_mx2_x2 1 1917 2 648 1594 35 mx2_x2
xsubckt_929_mx2_x2 1 1955 2 1624 116 1634 mx2_x2
xsubckt_928_mx2_x2 1 1956 2 1624 117 1642 mx2_x2
xsubckt_748_o2_x2 1 1774 2 1776 1784 o2_x2
xsubckt_1425_mx2_x2 1 1854 2 903 1229 52 mx2_x2
xsubckt_1826_sff1_x4 2 211 1 89 97 sff1_x4
xsubckt_1865_sff1_x4 2 202 1 1868 58 sff1_x4
xsubckt_1194_a2_x2 1 1428 2 284 577 a2_x2
xsubckt_1161_nand2_x0 2 1 1458 1459 700 nand2_x0
xsubckt_889_mx2_x2 1 1967 2 1662 144 1652 mx2_x2
xsubckt_888_mx2_x2 1 1652 2 563 1653 92 mx2_x2
xsubckt_694_nand3_x0 2 1 1825 262 269 132 nand3_x0
xsubckt_1382_mx2_x2 1 1858 2 903 1268 56 mx2_x2
xsubckt_1641_nand2_x0 2 1 1014 1015 1022 nand2_x0
xsubckt_1653_a2_x2 1 1002 2 1003 1005 a2_x2
xsubckt_1102_o2_x2 1 1503 2 1504 1527 o2_x2
xsubckt_906_nand3_x0 2 1 1638 889 895 158 nand3_x0
xsubckt_1478_a2_x2 1 1176 2 1177 1190 a2_x2
xsubckt_1673_a2_x2 1 982 2 983 985 a2_x2
xsubckt_1773_sff1_x4 2 208 1 1950 135 sff1_x4
xsubckt_867_nand2_x0 2 1 1670 1769 146 nand2_x0
xsubckt_297_nand2_x0 2 1 587 588 592 nand2_x0
xsubckt_30_inv_x0 2 1 111 883 inv_x0
xsubckt_31_inv_x0 2 1 13 882 inv_x0
xsubckt_32_inv_x0 2 1 66 881 inv_x0
xsubckt_33_inv_x0 2 1 68 880 inv_x0
xsubckt_160_nand2_x0 2 1 741 743 744 nand2_x0
xsubckt_1769_sff1_x4 2 205 1 179 28 sff1_x4
xcmpt_abc_11873_new_n335_hfns_3 2 1 905 901 buf_x4
xcmpt_abc_11873_new_n335_hfns_2 2 1 901 902 buf_x4
xcmpt_abc_11873_new_n335_hfns_1 2 1 901 903 buf_x4
xcmpt_abc_11873_new_n335_hfns_0 2 1 901 904 buf_x4
xsubckt_1103_nand2_x0 2 1 1502 1584 740 nand2_x0
xsubckt_798_ao22_x2 1 1729 2 1776 1784 148 ao22_x2
xsubckt_673_nand4_x0 2 1 218 220 221 222 223 nand4_x0
xsubckt_34_inv_x0 2 1 40 879 inv_x0
xsubckt_35_inv_x0 2 1 59 878 inv_x0
xsubckt_36_inv_x0 2 1 58 877 inv_x0
xsubckt_37_inv_x0 2 1 51 876 inv_x0
xsubckt_38_inv_x0 2 1 50 875 inv_x0
xsubckt_39_inv_x0 2 1 49 874 inv_x0
xsubckt_353_a4_x2 1 528 2 788 832 835 31 a4_x2
xsubckt_1276_nxr2_x1 1363 2 1 1365 1373 nxr2_x1
xsubckt_1191_nand2_x0 2 1 1431 1435 1437 nand2_x0
xsubckt_198_a4_x2 1 693 2 694 700 704 709 a4_x2
xsubckt_433_oa22_x2 1 449 2 713 497 554 oa22_x2
xsubckt_456_nand3_x0 2 1 426 680 703 718 nand3_x0
xsubckt_632_ao22_x2 1 256 2 710 565 484 ao22_x2
xsubckt_1528_ao22_x2 1 1127 2 1141 1143 1189 ao22_x2
xsubckt_1567_ao22_x2 1 1088 2 891 1202 1089 ao22_x2
xsubckt_1725_oa22_x2 1 930 2 931 1144 1157 oa22_x2
xsubckt_1169_nor3_x0 2 1 1451 106 159 36 nor3_x0
xsubckt_1009_nand3_x0 2 1 1576 1577 1578 650 nand3_x0
xsubckt_846_nand3_x0 2 1 1688 1767 1775 55 nand3_x0
xsubckt_760_nand2_x0 2 1 1762 1763 1764 nand2_x0
xsubckt_190_nand2_x0 2 1 704 707 713 nand2_x0
xsubckt_324_a2_x2 1 560 2 561 567 a2_x2
xsubckt_461_a3_x2 2 421 1 698 792 799 a3_x2
xsubckt_471_a3_x2 2 411 1 412 422 429 a3_x2
xsubckt_1530_nand3_x0 2 1 1125 1140 1142 1176 nand3_x0
xsubckt_970_a3_x2 2 1609 1 628 731 734 a3_x2
xsubckt_756_nand3_x0 2 1 1766 1767 1775 59 nand3_x0
xsubckt_149_a2_x2 1 755 2 757 759 a2_x2
xsubckt_159_a2_x2 1 742 2 743 744 a2_x2
xsubckt_344_a2_x2 1 537 2 543 713 a2_x2
xsubckt_364_a2_x2 1 517 2 518 520 a2_x2
xsubckt_1350_nand3_x0 2 1 1297 773 780 175 nand3_x0
xsubckt_1051_a4_x2 1 1544 2 650 742 747 761 a4_x2
xsubckt_873_a2_x2 1 1666 2 1668 67 a2_x2
xsubckt_1309_nand3_x0 2 1 1334 773 780 163 nand3_x0
xsubckt_1650_nand3_x0 2 1 1005 698 795 58 nand3_x0
xsubckt_1248_a3_x2 2 1390 1 471 553 594 a3_x2
xsubckt_839_nand2_x0 2 1 1982 1694 1698 nand2_x0
xsubckt_790_nand2_x0 2 1 1736 1774 149 nand2_x0
xsubckt_768_oa22_x2 1 1755 2 536 657 808 oa22_x2
xsubckt_641_oa22_x2 1 247 2 249 550 883 oa22_x2
xsubckt_218_nand3_x0 2 1 669 681 712 724 nand3_x0
xsubckt_396_nand3_x0 2 1 485 497 681 794 nand3_x0
xsubckt_1433_nand2_x0 2 1 1221 672 106 nand2_x0
xsubckt_1519_nand3_x0 2 1 1136 1138 1139 1160 nand3_x0
xsubckt_1811_sff1_x4 2 209 1 1913 159 sff1_x4
xsubckt_1850_sff1_x4 2 202 1 1883 166 sff1_x4
xsubckt_1233_mx2_x2 1 1881 2 1394 1974 164 mx2_x2
xsubckt_1232_mx2_x2 1 1882 2 1394 1975 165 mx2_x2
xsubckt_1231_mx2_x2 1 1883 2 1394 1976 166 mx2_x2
xsubckt_1230_mx2_x2 1 1884 2 1394 1983 167 mx2_x2
xsubckt_1052_a2_x2 1 1543 2 1609 621 a2_x2
xsubckt_686_o2_x2 1 1832 2 256 860 o2_x2
xsubckt_125_nor2_x0 2 1 785 25 31 nor2_x0
xsubckt_1473_a3_x2 2 1181 1 1182 1183 1185 a3_x2
xsubckt_1807_sff1_x4 2 205 1 1917 35 sff1_x4
xsubckt_1846_sff1_x4 2 209 1 1841 158 sff1_x4
xsubckt_1885_sff1_x4 2 202 1 1848 150 sff1_x4
xsubckt_1239_mx2_x2 1 1875 2 1394 1982 174 mx2_x2
xsubckt_1238_mx2_x2 1 1876 2 1394 1969 175 mx2_x2
xsubckt_1237_mx2_x2 1 1877 2 1394 1970 176 mx2_x2
xsubckt_1236_mx2_x2 1 1878 2 1394 1971 161 mx2_x2
xsubckt_1235_mx2_x2 1 1879 2 1394 1972 162 mx2_x2
xsubckt_1234_mx2_x2 1 1880 2 1394 1973 163 mx2_x2
xsubckt_1158_o4_x2 1 1461 2 1466 1667 112 106 o4_x2
xsubckt_1092_a2_x2 1 1905 2 1511 1516 a2_x2
xsubckt_696_nand3_x0 2 1 1823 262 268 116 nand3_x0
xsubckt_676_oa22_x2 1 215 2 253 700 892 oa22_x2
xsubckt_518_nand3_x0 2 1 365 570 718 800 nand3_x0
xsubckt_569_nor3_x0 2 1 315 399 482 490 nor3_x0
xsubckt_1339_nand3_x0 2 1 1307 773 780 176 nand3_x0
xsubckt_1445_oa22_x2 1 1209 2 718 707 528 oa22_x2
xsubckt_1541_a2_x2 1 1114 2 1115 1117 a2_x2
xsubckt_1628_mx2_x2 1 1027 2 1030 1176 1189 mx2_x2
xsubckt_201_nand3_x0 2 1 690 691 708 831 nand3_x0
xsubckt_506_nxr2_x1 377 2 1 742 747 nxr2_x1
xsubckt_1754_sff1_x4 2 207 1 1963 140 sff1_x4
xsubckt_1793_sff1_x4 2 209 1 1931 43 sff1_x4
xsubckt_822_nand2_x0 2 1 1708 1780 93 nand2_x0
xsubckt_1789_sff1_x4 2 211 1 1935 105 sff1_x4
xsubckt_1710_nxr2_x1 945 2 1 953 956 nxr2_x1
xsubckt_162_nand2_x0 2 1 739 741 749 nand2_x0
xsubckt_299_nand2_x0 2 1 585 597 718 nand2_x0
xsubckt_869_nand2_x0 2 1 1977 1669 1673 nand2_x0
xcmpt_abc_11873_new_n532_hfns_3 2 1 682 678 buf_x4
xcmpt_abc_11873_new_n532_hfns_2 2 1 678 679 buf_x4
xcmpt_abc_11873_new_n532_hfns_1 2 1 678 680 buf_x4
xcmpt_abc_11873_new_n532_hfns_0 2 1 678 681 buf_x4
xsubckt_552_nand2_x0 2 1 332 522 800 nand2_x0
xsubckt_271_a4_x2 1 613 2 620 628 729 766 a4_x2
xfeed_19 2 1 decap_w0
xfeed_18 2 1 decap_w0
xfeed_17 2 1 decap_w0
xfeed_16 2 1 decap_w0
xfeed_15 2 1 decap_w0
xfeed_14 2 1 decap_w0
xfeed_13 2 1 decap_w0
xfeed_12 2 1 decap_w0
xfeed_11 2 1 decap_w0
xfeed_10 2 1 decap_w0
xsubckt_1460_ao22_x2 1 1194 2 1800 1206 1196 ao22_x2
xsubckt_1025_ao22_x2 1 1920 2 1574 1569 1563 ao22_x2
xsubckt_1193_nor3_x0 2 1 1429 1431 1432 1439 nor3_x0
xsubckt_1279_nand3_x0 2 1 1361 773 780 166 nand3_x0
xsubckt_623_a3_x2 2 265 1 266 276 282 a3_x2
xsubckt_595_a4_x2 1 291 2 292 295 338 531 a4_x2
xsubckt_428_a3_x2 2 454 1 456 729 766 a3_x2
xsubckt_762_nand2_x0 2 1 1760 1761 1766 nand2_x0
xfeed_29 2 1 decap_w0
xfeed_28 2 1 decap_w0
xfeed_27 2 1 decap_w0
xfeed_26 2 1 tie
xfeed_25 2 1 decap_w0
xfeed_24 2 1 decap_w0
xfeed_23 2 1 decap_w0
xfeed_22 2 1 decap_w0
xfeed_21 2 1 decap_w0
xfeed_20 2 1 decap_w0
xsubckt_1456_ao22_x2 1 1198 2 802 1200 1233 ao22_x2
xsubckt_1352_nand3_x0 2 1 1295 591 792 175 nand3_x0
xsubckt_272_a2_x2 1 612 2 741 747 a2_x2
xsubckt_576_a2_x2 1 309 2 322 458 a2_x2
xsubckt_556_a2_x2 1 328 2 329 331 a2_x2
xsubckt_492_nand2_x0 2 1 182 391 410 nand2_x0
xsubckt_188_nand3_x0 2 1 706 708 26 836 nand3_x0
xsubckt_668_nand3_x0 2 1 223 262 268 118 nand3_x0
xsubckt_751_a2_x2 1 1771 2 1773 700 a2_x2
xsubckt_792_oa22_x2 1 1734 2 536 657 805 oa22_x2
xsubckt_987_a3_x2 2 1597 1 461 612 761 a3_x2
xfeed_39 2 1 decap_w0
xfeed_38 2 1 tie
xfeed_37 2 1 tie
xfeed_36 2 1 decap_w0
xfeed_35 2 1 decap_w0
xfeed_34 2 1 decap_w0
xfeed_33 2 1 decap_w0
xfeed_32 2 1 decap_w0
xfeed_31 2 1 decap_w0
xfeed_30 2 1 decap_w0
xsubckt_1652_nand3_x0 2 1 1003 1181 1186 92 nand3_x0
xsubckt_1615_nand2_x0 2 1 1040 1041 1286 nand2_x0
xsubckt_1525_nand2_x0 2 1 1130 1132 1133 nand2_x0
xsubckt_1522_oa22_x2 1 1133 2 1204 1790 888 oa22_x2
xsubckt_210_o2_x2 1 677 2 4 9 o2_x2
xsubckt_714_oa22_x2 1 1806 2 249 550 882 oa22_x2
xsubckt_972_nand2_x0 2 1 1928 1608 1610 nand2_x0
xsubckt_1038_a4_x2 1 1554 2 783 795 20 9 a4_x2
xsubckt_1045_nand2_x0 2 1 1915 1548 1552 nand2_x0
xsubckt_1172_nand3_x0 2 1 1448 703 719 36 nand3_x0
xsubckt_1253_a4_x2 1 1385 2 1783 577 593 709 a4_x2
xsubckt_1870_sff1_x4 2 202 1 1863 47 sff1_x4
xsubckt_1831_sff1_x4 2 209 1 1901 72 sff1_x4
xsubckt_1721_ao22_x2 1 934 2 936 937 1092 ao22_x2
xsubckt_1489_nor3_x0 2 1 1165 1167 1168 289 nor3_x0
xsubckt_1435_nand2_x0 2 1 1219 1220 1772 nand2_x0
xsubckt_930_mx2_x2 1 1954 2 1624 115 1629 mx2_x2
xsubckt_931_mx2_x2 1 1953 2 1624 114 1625 mx2_x2
xsubckt_933_mx2_x2 1 1952 2 1623 137 1661 mx2_x2
xsubckt_934_mx2_x2 1 1951 2 1623 136 1652 mx2_x2
xsubckt_1168_nand4_x0 2 1 1452 784 788 794 911 nand4_x0
xfeed_46 2 1 decap_w0
xfeed_45 2 1 decap_w0
xfeed_44 2 1 decap_w0
xfeed_43 2 1 decap_w0
xfeed_42 2 1 decap_w0
xfeed_41 2 1 decap_w0
xfeed_40 2 1 decap_w0
xsubckt_1866_sff1_x4 2 202 1 1867 51 sff1_x4
xsubckt_1562_mx3_x2 2 1 1093 1226 1101 1129 1096 1099 mx3_x2
xsubckt_1561_mx3_x2 2 1 1094 1226 1101 1128 1095 1100 mx3_x2
xsubckt_1345_nand2_x0 2 1 1301 1303 1309 nand2_x0
xsubckt_561_nand3_x0 2 1 323 437 454 645 nand3_x0
xsubckt_401_nor4_x0 2 1 480 23 19 26 31 nor4_x0
xsubckt_935_mx2_x2 1 1950 2 1623 135 1647 mx2_x2
xsubckt_936_mx2_x2 1 1949 2 1623 134 1643 mx2_x2
xsubckt_937_mx2_x2 1 1948 2 1623 133 1642 mx2_x2
xsubckt_938_mx2_x2 1 1947 2 1623 132 1634 mx2_x2
xsubckt_939_mx2_x2 1 1946 2 1623 131 1629 mx2_x2
xsubckt_1196_a3_x2 2 1426 1 583 589 700 a3_x2
xfeed_49 2 1 decap_w0
xfeed_48 2 1 decap_w0
xfeed_47 2 1 decap_w0
xsubckt_1827_sff1_x4 2 211 1 88 96 sff1_x4
xsubckt_434_nand2_x0 2 1 448 640 693 nand2_x0
xsubckt_894_mx2_x2 1 1647 2 563 1648 91 mx2_x2
xsubckt_895_mx2_x2 1 1966 2 1662 143 1647 mx2_x2
xsubckt_1114_nand3_x0 2 1 1901 1493 398 518 nand3_x0
xsubckt_1151_nand4_x0 2 1 1467 1492 585 700 777 nand4_x0
xsubckt_1175_mx3_x2 2 1 1445 1451 42 155 153 910 mx3_x2
xsubckt_1274_a2_x2 1 1365 2 1366 1370 a2_x2
xfeed_53 2 1 decap_w0
xfeed_52 2 1 decap_w0
xfeed_51 2 1 decap_w0
xfeed_50 2 1 decap_w0
xsubckt_1774_sff1_x4 2 208 1 1949 134 sff1_x4
xsubckt_1392_mx2_x2 1 1857 2 903 1259 55 mx2_x2
xsubckt_381_nand3_x0 2 1 500 610 612 767 nand3_x0
xsubckt_824_nand2_x0 2 1 1706 1707 176 nand2_x0
xsubckt_899_mx2_x2 1 1643 2 563 1644 90 mx2_x2
xsubckt_1048_mx2_x2 1 1913 2 1553 1551 159 mx2_x2
xfeed_59 2 1 decap_w0
xfeed_58 2 1 tie
xfeed_57 2 1 decap_w0
xfeed_56 2 1 decap_w0
xfeed_55 2 1 decap_w0
xfeed_54 2 1 decap_w0
xsubckt_1730_nxr2_x1 925 2 1 932 934 nxr2_x1
xsubckt_1699_ao22_x2 1 956 2 959 961 987 ao22_x2
xsubckt_1334_oa22_x2 1 1311 2 1327 1319 1314 oa22_x2
xsubckt_40_inv_x0 2 1 48 873 inv_x0
xsubckt_241_ao22_x2 1 643 2 772 768 645 ao22_x2
xsubckt_681_nand3_x0 2 1 1837 262 268 117 nand3_x0
xfeed_60 2 1 decap_w0
xsubckt_1726_nxr2_x1 929 2 1 930 1145 nxr2_x1
xsubckt_1506_o2_x2 1 1149 2 1200 809 o2_x2
xsubckt_41_inv_x0 2 1 47 872 inv_x0
xsubckt_42_inv_x0 2 1 46 871 inv_x0
xsubckt_43_inv_x0 2 1 63 870 inv_x0
xsubckt_44_inv_x0 2 1 62 869 inv_x0
xsubckt_45_inv_x0 2 1 61 868 inv_x0
xsubckt_46_inv_x0 2 1 60 867 inv_x0
xsubckt_1266_nor3_x0 2 1 1372 1374 1376 1388 nor3_x0
xfeed_69 2 1 decap_w0
xfeed_68 2 1 decap_w0
xfeed_67 2 1 decap_w0
xfeed_66 2 1 decap_w0
xfeed_65 2 1 decap_w0
xfeed_64 2 1 decap_w0
xfeed_63 2 1 tie
xfeed_62 2 1 decap_w0
xfeed_61 2 1 decap_w0
xsubckt_1675_nand2_x0 2 1 980 981 1160 nand2_x0
xsubckt_1568_ao22_x2 1 1087 2 1834 1206 1088 ao22_x2
xsubckt_1369_oa22_x2 1 1279 2 1300 1291 1282 oa22_x2
xsubckt_409_nand4_x0 2 1 472 473 476 477 481 nand4_x0
xsubckt_374_nand2_x0 2 1 507 707 718 nand2_x0
xsubckt_323_nand3_x0 2 1 561 566 713 800 nand3_x0
xsubckt_47_inv_x0 2 1 43 866 inv_x0
xsubckt_48_inv_x0 2 1 45 865 inv_x0
xsubckt_49_inv_x0 2 1 44 864 inv_x0
xsubckt_1054_nand3_x0 2 1 1912 1542 1545 1546 nand3_x0
xsubckt_1645_nor2_x0 2 1 1010 1011 1013 nor2_x0
xsubckt_1585_nand2_x0 2 1 1070 1071 1154 nand2_x0
xsubckt_571_a3_x2 2 313 1 318 422 429 a3_x2
xsubckt_541_a3_x2 2 342 1 343 498 571 a3_x2
xsubckt_521_a3_x2 2 362 1 363 364 365 a3_x2
xsubckt_376_a3_x2 2 505 1 612 617 753 a3_x2
xsubckt_120_a2_x2 1 801 2 900 9 a2_x2
xsubckt_233_nand3_x0 2 1 654 656 657 663 nand3_x0
xsubckt_319_nand4_x0 2 1 565 833 20 835 31 nand4_x0
xsubckt_764_nand2_x0 2 1 1759 1792 240 nand2_x0
xsubckt_854_nand2_x0 2 1 1681 1769 148 nand2_x0
xfeed_79 2 1 decap_w0
xfeed_78 2 1 decap_w0
xfeed_77 2 1 decap_w0
xfeed_76 2 1 decap_w0
xfeed_75 2 1 tie
xfeed_74 2 1 decap_w0
xfeed_73 2 1 tie
xfeed_72 2 1 decap_w0
xfeed_71 2 1 decap_w0
xfeed_70 2 1 decap_w0
xsubckt_591_a3_x2 2 295 1 296 297 298 a3_x2
xsubckt_581_a3_x2 2 304 1 305 306 344 a3_x2
xsubckt_180_nand4_x0 2 1 721 788 831 26 836 nand4_x0
xsubckt_194_nand2_x0 2 1 700 703 719 nand2_x0
xsubckt_239_a2_x2 1 645 2 650 900 a2_x2
xsubckt_1707_nand2_x0 2 1 948 672 160 nand2_x0
xsubckt_1542_nxr2_x1 1113 2 1 1114 1164 nxr2_x1
xsubckt_443_nand3_x0 2 1 439 591 681 712 nand3_x0
xsubckt_406_nand2_x0 2 1 475 480 832 nand2_x0
xsubckt_279_a2_x2 1 605 2 606 631 a2_x2
xsubckt_316_nand2_x0 2 1 568 570 712 nand2_x0
xsubckt_913_a2_x2 1 1632 2 1640 888 a2_x2
xfeed_89 2 1 decap_w0
xfeed_88 2 1 decap_w0
xfeed_87 2 1 decap_w0
xfeed_86 2 1 decap_w0
xfeed_85 2 1 decap_w0
xfeed_84 2 1 decap_w0
xfeed_83 2 1 decap_w0
xfeed_82 2 1 decap_w0
xfeed_81 2 1 decap_w0
xfeed_80 2 1 decap_w0
xsubckt_1503_oa22_x2 1 1853 2 1152 1156 1228 oa22_x2
xsubckt_1448_nor4_x0 2 1 1206 1207 1208 1421 281 nor4_x0
xsubckt_207_o2_x2 1 684 2 14 155 o2_x2
xsubckt_212_nand4_x0 2 1 675 784 787 831 27 nand4_x0
xsubckt_226_nand2_x0 2 1 661 17 27 nand2_x0
xsubckt_773_oa22_x2 1 1751 2 1770 1771 854 oa22_x2
xsubckt_1084_nand3_x0 2 1 1517 1518 1528 1583 nand3_x0
xsubckt_1181_a4_x2 1 1441 2 784 832 23 834 a4_x2
xsubckt_1890_sff1_x4 2 202 1 1843 154 sff1_x4
xsubckt_1851_sff1_x4 2 206 1 1882 165 sff1_x4
xsubckt_1812_sff1_x4 2 209 1 1912 82 sff1_x4
xsubckt_1474_nand3_x0 2 1 1180 1181 1186 86 nand3_x0
xsubckt_412_o2_x2 1 469 2 663 677 o2_x2
xfeed_99 2 1 tie
xfeed_98 2 1 decap_w0
xfeed_97 2 1 decap_w0
xfeed_96 2 1 tie
xfeed_95 2 1 decap_w0
xfeed_94 2 1 decap_w0
xfeed_93 2 1 tie
xfeed_92 2 1 tie
xfeed_91 2 1 tie
xfeed_90 2 1 decap_w0
xsubckt_1886_sff1_x4 2 202 1 1847 149 sff1_x4
xsubckt_1632_mx2_x2 1 1023 2 1037 1025 1029 mx2_x2
xsubckt_1631_mx2_x2 1 1024 2 1037 1026 1028 mx2_x2
xsubckt_1384_nand3_x0 2 1 1266 773 780 172 nand3_x0
xsubckt_165_nor2_x0 2 1 736 86 71 nor2_x0
xsubckt_690_nand4_x0 2 1 1828 1829 1830 1832 249 nand4_x0
xsubckt_726_o2_x2 1 1795 2 256 857 o2_x2
xsubckt_1112_a2_x2 1 1494 2 900 71 a2_x2
xsubckt_1132_a2_x2 1 1483 2 147 42 a2_x2
xsubckt_1240_mx2_x2 1 1874 2 1394 1981 173 mx2_x2
xsubckt_1257_nand2_x0 2 1 1381 1383 777 nand2_x0
xsubckt_1847_sff1_x4 2 210 1 1886 113 sff1_x4
xsubckt_1808_sff1_x4 2 209 1 1916 106 sff1_x4
xsubckt_1634_mx2_x2 1 1021 2 1227 1024 1063 mx2_x2
xsubckt_1633_mx2_x2 1 1022 2 1227 1023 1062 mx2_x2
xsubckt_1426_a2_x2 1 1228 2 156 903 a2_x2
xsubckt_638_oa22_x2 1 250 2 253 700 897 oa22_x2
xsubckt_473_nand3_x0 2 1 409 543 680 713 nand3_x0
xsubckt_436_nand2_x0 2 1 446 543 718 nand2_x0
xsubckt_422_nand4_x0 2 1 460 621 627 729 766 nand4_x0
xsubckt_649_nand4_x0 2 1 240 242 243 244 245 nand4_x0
xsubckt_677_oa22_x2 1 1840 2 249 550 914 oa22_x2
xsubckt_1241_mx2_x2 1 1873 2 1394 1980 172 mx2_x2
xsubckt_1242_mx2_x2 1 1872 2 1394 1979 171 mx2_x2
xsubckt_1243_mx2_x2 1 1871 2 1394 1978 170 mx2_x2
xsubckt_1244_mx2_x2 1 1870 2 1394 1977 169 mx2_x2
xsubckt_1794_sff1_x4 2 210 1 1930 110 sff1_x4
xsubckt_1755_sff1_x4 2 207 1 1962 139 sff1_x4
xsubckt_1691_a2_x2 1 964 2 971 980 a2_x2
xsubckt_1681_a2_x2 1 974 2 975 1174 a2_x2
xsubckt_722_nand4_x0 2 1 1799 1801 1802 1803 1804 nand4_x0
xsubckt_1711_nxr2_x1 944 2 1 953 955 nxr2_x1
xsubckt_1599_mx2_x2 1 1056 2 1058 1176 1189 mx2_x2
xsubckt_1594_nand3_x0 2 1 1061 698 792 50 nand3_x0
xsubckt_683_nand3_x0 2 1 1835 262 269 133 nand3_x0
xsubckt_1630_nand2_x0 2 1 1025 1027 1174 nand2_x0
xsubckt_1592_ao22_x2 1 1063 2 219 1206 1065 ao22_x2
xsubckt_1553_ao22_x2 1 1102 2 1821 1206 1104 ao22_x2
xsubckt_1315_oa22_x2 1 1328 2 48 1377 1330 oa22_x2
xsubckt_199_nand4_x0 2 1 692 694 700 704 709 nand4_x0
xsubckt_1588_ao22_x2 1 1067 2 806 1200 1274 ao22_x2
xsubckt_1549_ao22_x2 1 1106 2 804 1200 1255 ao22_x2
xsubckt_1297_nxr2_x1 1344 2 1 1347 1355 nxr2_x1
xsubckt_452_nand4_x0 2 1 430 462 612 645 753 nand4_x0
xsubckt_1422_ao22_x2 1 1231 2 802 1387 1232 ao22_x2
xsubckt_1360_nand2_x0 2 1 1288 1386 91 nand2_x0
xsubckt_130_ao22_x2 1 774 2 83 861 913 ao22_x2
xsubckt_244_a3_x2 2 640 1 655 659 800 a3_x2
xsubckt_766_nand2_x0 2 1 1757 1774 152 nand2_x0
xsubckt_818_nor2_x0 2 1 1711 1712 1715 nor2_x0
xsubckt_890_a4_x2 1 1651 2 151 154 160 158 a4_x2
xsubckt_606_a2_x2 1 282 2 283 633 a2_x2
xsubckt_147_a2_x2 1 757 2 758 774 a2_x2
xsubckt_137_a2_x2 1 767 2 770 776 a2_x2
xsubckt_688_ao22_x2 1 1830 2 891 252 1831 ao22_x2
xsubckt_408_nand2_x0 2 1 473 474 800 nand2_x0
xsubckt_1139_nand2_x0 2 1 1477 1478 444 nand2_x0
xsubckt_976_nand2_x0 2 1 1605 648 108 nand2_x0
xsubckt_1871_sff1_x4 2 202 1 1862 46 sff1_x4
xsubckt_1832_sff1_x4 2 211 1 1900 80 sff1_x4
xsubckt_1401_a3_x2 2 1250 1 1251 1260 1269 a3_x2
xsubckt_1390_nand2_x0 2 1 1260 1262 1267 nand2_x0
xsubckt_1353_a4_x2 1 1294 2 1295 1296 1297 550 a4_x2
xsubckt_145_o2_x2 1 759 2 90 71 o2_x2
xsubckt_138_nand2_x0 2 1 766 770 776 nand2_x0
xsubckt_872_nand4_x0 2 1 1667 784 788 794 909 nand4_x0
xsubckt_940_mx2_x2 1 1945 2 1623 130 1625 mx2_x2
xsubckt_1000_a2_x2 1 1585 2 620 730 a2_x2
xsubckt_1010_a2_x2 1 1575 2 1600 620 a2_x2
xspare_buffer_9 2 1 212 207 buf_x4
xspare_buffer_8 2 1 212 208 buf_x4
xspare_buffer_7 2 1 7 6 buf_x4
xspare_buffer_6 2 1 212 209 buf_x4
xspare_buffer_5 2 1 212 210 buf_x4
xspare_buffer_4 2 1 212 211 buf_x4
xspare_buffer_3 2 1 8 7 buf_x4
xspare_buffer_0 2 1 213 212 buf_x4
xsubckt_1471_a3_x2 2 1183 1 1184 284 577 a3_x2
xsubckt_1441_a3_x2 2 1213 1 1215 1216 1217 a3_x2
xsubckt_1349_nand2_x0 2 1 1298 1379 44 nand2_x0
xsubckt_301_nand2_x0 2 1 583 591 717 nand2_x0
xsubckt_662_oa22_x2 1 228 2 486 568 876 oa22_x2
xsubckt_942_mx2_x2 1 1944 2 1622 129 1661 mx2_x2
xsubckt_943_mx2_x2 1 1943 2 1622 128 1652 mx2_x2
xsubckt_944_mx2_x2 1 1942 2 1622 127 1647 mx2_x2
xsubckt_945_mx2_x2 1 1941 2 1622 126 1643 mx2_x2
xsubckt_946_mx2_x2 1 1940 2 1622 125 1642 mx2_x2
xsubckt_947_mx2_x2 1 1939 2 1622 124 1634 mx2_x2
xsubckt_1273_ao22_x2 1 1366 2 896 1385 1367 ao22_x2
xsubckt_1867_sff1_x4 2 202 1 1866 50 sff1_x4
xsubckt_1828_sff1_x4 2 211 1 87 95 sff1_x4
xsubckt_1718_ao22_x2 1 937 2 940 941 1069 ao22_x2
xsubckt_1690_nand2_x0 2 1 965 967 1212 nand2_x0
xsubckt_1344_a2_x2 1 1302 2 1303 1309 a2_x2
xsubckt_441_nor4_x0 2 1 441 442 443 447 672 nor4_x0
xsubckt_438_nand2_x0 2 1 444 688 718 nand2_x0
xsubckt_948_mx2_x2 1 1938 2 1622 123 1629 mx2_x2
xsubckt_949_mx2_x2 1 1937 2 1622 122 1625 mx2_x2
xsubckt_1032_nand2_x0 2 1 1918 1560 1562 nand2_x0
xsubckt_1159_a2_x2 1 1460 2 1461 1468 a2_x2
xsubckt_1658_a2_x2 1 997 2 998 1174 a2_x2
xsubckt_1626_ao22_x2 1 1029 2 1033 1035 1189 ao22_x2
xsubckt_121_nand2_x0 2 1 797 900 9 nand2_x0
xsubckt_992_nand4_x0 2 1 1593 628 729 742 747 nand4_x0
xsubckt_1056_mx2_x2 1 1911 2 648 1541 68 mx2_x2
xsubckt_1189_a2_x2 1 1433 2 541 667 a2_x2
xsubckt_1775_sff1_x4 2 208 1 1948 133 sff1_x4
xsubckt_1418_nand3_x0 2 1 1235 773 780 169 nand3_x0
xsubckt_1328_nand3_x0 2 1 1317 773 780 161 nand3_x0
xsubckt_1379_nand2_x0 2 1 1270 1272 1277 nand2_x0
xsubckt_50_inv_x0 2 1 57 863 inv_x0
xsubckt_51_inv_x0 2 1 56 862 inv_x0
xsubckt_52_inv_x0 2 1 177 861 inv_x0
xsubckt_53_inv_x0 2 1 55 860 inv_x0
xsubckt_1192_nor4_x0 2 1 1430 1434 1436 1440 1441 nor4_x0
xsubckt_1646_o2_x2 1 1009 2 1011 1013 o2_x2
xsubckt_454_nand4_x0 2 1 428 741 749 754 760 nand4_x0
xsubckt_54_inv_x0 2 1 54 859 inv_x0
xsubckt_55_inv_x0 2 1 53 858 inv_x0
xsubckt_56_inv_x0 2 1 52 857 inv_x0
xsubckt_57_inv_x0 2 1 168 856 inv_x0
xsubckt_58_inv_x0 2 1 167 855 inv_x0
xsubckt_59_inv_x0 2 1 166 854 inv_x0
xsubckt_318_a4_x2 1 566 2 833 19 835 31 a4_x2
xsubckt_919_nxr2_x1 1627 2 1 1639 887 nxr2_x1
xsubckt_985_nand3_x0 2 1 1598 1600 1614 621 nand3_x0
xsubckt_1062_nand2_x0 2 1 1909 1537 1539 nand2_x0
xsubckt_1185_nand4_x0 2 1 1437 784 831 27 23 nand4_x0
xsubckt_1674_nxr2_x1 981 2 1 982 1164 nxr2_x1
xsubckt_1589_nand2_x0 2 1 1066 1068 1274 nand2_x0
xsubckt_1538_nand3_x0 2 1 1117 697 795 48 nand3_x0
xsubckt_426_a3_x2 2 456 1 623 625 628 a3_x2
xsubckt_200_a2_x2 1 691 2 26 31 a2_x2
xsubckt_717_nand3_x0 2 1 1804 263 268 122 nand3_x0
xsubckt_1204_oa22_x2 1 1418 2 496 695 790 oa22_x2
xspare_feed_13 2 1 decap_w0
xspare_feed_12 2 1 decap_w0
xspare_feed_11 2 1 decap_w0
xspare_feed_10 2 1 decap_w0
xsubckt_1635_nxr2_x1 1020 2 1 1031 1164 nxr2_x1
xsubckt_627_nand3_x0 2 1 261 262 269 137 nand3_x0
xsubckt_524_a2_x2 1 359 2 360 361 a2_x2
xsubckt_329_a2_x2 1 555 2 556 558 a2_x2
xsubckt_905_a3_x2 2 1639 1 889 895 158 a3_x2
xsubckt_1221_nand3_x0 2 1 1401 1404 279 539 nand3_x0
xsubckt_1278_oa22_x2 1 1362 2 1380 579 876 oa22_x2
xspare_feed_19 2 1 decap_w0
xspare_feed_18 2 1 decap_w0
xspare_feed_17 2 1 decap_w0
xspare_feed_16 2 1 decap_w0
xspare_feed_15 2 1 decap_w0
xspare_feed_14 2 1 decap_w0
xsubckt_785_nor2_x0 2 1 1740 1741 1744 nor2_x0
xsubckt_841_nand2_x0 2 1 1692 1707 173 nand2_x0
xsubckt_1217_nand4_x0 2 1 1405 1406 1407 671 690 nand4_x0
xspare_feed_20 2 1 decap_w0
xsubckt_1543_nxr2_x1 1112 2 1 1114 1165 nxr2_x1
xsubckt_1431_nand3_x0 2 1 1223 672 880 912 nand3_x0
xsubckt_498_nand2_x0 2 1 385 453 616 nand2_x0
xsubckt_216_nand4_x0 2 1 671 788 794 26 836 nand4_x0
xsubckt_774_oa22_x2 1 1750 2 536 657 807 oa22_x2
xsubckt_978_nand2_x0 2 1 1926 1604 1605 nand2_x0
xspare_feed_25 2 1 tie
xspare_feed_24 2 1 tie
xspare_feed_23 2 1 decap_w0
xspare_feed_22 2 1 tie
xspare_feed_21 2 1 tie
xsubckt_1891_sff1_x4 2 202 1 1842 157 sff1_x4
xsubckt_1703_ao22_x2 1 952 2 954 956 1014 ao22_x2
xsubckt_532_o2_x2 1 351 2 656 677 o2_x2
xsubckt_258_nor2_x0 2 1 626 88 71 nor2_x0
xsubckt_875_o4_x2 1 1664 2 1665 1666 278 563 o4_x2
xsubckt_1020_oa22_x2 1 1566 2 740 615 378 oa22_x2
xsubckt_1088_nand3_x0 2 1 1514 1515 1541 612 nand3_x0
xsubckt_1096_a4_x2 1 1507 2 1508 1509 1514 1583 a4_x2
xsubckt_1214_nand2_x0 2 1 1408 1409 709 nand2_x0
xspare_feed_9 2 1 decap_w0
xspare_feed_8 2 1 decap_w0
xspare_feed_7 2 1 decap_w0
xspare_feed_6 2 1 decap_w0
xspare_feed_5 2 1 decap_w0
xspare_feed_4 2 1 decap_w0
xspare_feed_3 2 1 decap_w0
xspare_feed_2 2 1 decap_w0
xspare_feed_1 2 1 decap_w0
xspare_feed_0 2 1 decap_w0
xsubckt_1852_sff1_x4 2 207 1 1881 164 sff1_x4
xsubckt_1813_sff1_x4 2 209 1 1911 68 sff1_x4
xsubckt_1438_a3_x2 2 1216 1 1404 519 583 a3_x2
xsubckt_357_o2_x2 1 524 2 525 797 o2_x2
xsubckt_643_oa22_x2 1 191 2 288 257 246 oa22_x2
xsubckt_657_nand3_x0 2 1 233 263 269 143 nand3_x0
xsubckt_1037_a2_x2 1 1916 2 1555 1557 a2_x2
xsubckt_1887_sff1_x4 2 202 1 1846 148 sff1_x4
xsubckt_1848_sff1_x4 2 202 1 1885 168 sff1_x4
xsubckt_1809_sff1_x4 2 209 1 1915 160 sff1_x4
xsubckt_1760_sff1_x4 2 207 1 1957 118 sff1_x4
xsubckt_1701_a2_x2 1 954 2 1017 1021 a2_x2
xsubckt_1692_nand2_x0 2 1 963 971 980 nand2_x0
xsubckt_1282_a2_x2 1 1358 2 1359 1361 a2_x2
xsubckt_391_nand2_x0 2 1 490 491 495 nand2_x0
xsubckt_1034_nand2_x0 2 1 1557 648 906 nand2_x0
xsubckt_1057_a2_x2 1 1540 2 648 12 a2_x2
xsubckt_1077_a2_x2 1 1907 2 1524 1533 a2_x2
xsubckt_1097_a2_x2 1 1506 2 1507 1520 a2_x2
xsubckt_1272_a2_x2 1 1367 2 1368 1369 a2_x2
xsubckt_603_nand2_x0 2 1 0 285 288 nand2_x0
xsubckt_730_nand3_x0 2 1 1792 283 290 633 nand3_x0
xsubckt_1795_sff1_x4 2 211 1 1929 39 sff1_x4
xsubckt_1756_sff1_x4 2 208 1 1961 138 sff1_x4
xsubckt_1607_ao22_x2 1 1048 2 1161 1051 1154 ao22_x2
xsubckt_1596_a2_x2 1 1059 2 1060 1061 a2_x2
xsubckt_1226_nor4_x0 2 1 1396 1397 1403 1405 1408 nor4_x0
xsubckt_1504_o2_x2 1 1151 2 155 9 o2_x2
xsubckt_1281_nand3_x0 2 1 1359 1360 566 793 nand3_x0
xsubckt_421_a4_x2 1 461 2 621 627 729 766 a4_x2
xsubckt_419_nand3_x0 2 1 463 566 680 712 nand3_x0
xsubckt_333_nand2_x0 2 1 551 566 793 nand2_x0
xsubckt_687_nand3_x0 2 1 1831 566 775 793 nand3_x0
xsubckt_1197_ao22_x2 1 1425 2 718 712 543 ao22_x2
xsubckt_1712_oa22_x2 1 943 2 944 946 948 oa22_x2
xsubckt_1708_nxr2_x1 947 2 1 957 960 nxr2_x1
xsubckt_276_a4_x2 1 608 2 741 747 754 760 a4_x2
xsubckt_1031_ao22_x2 1 1558 2 761 755 650 ao22_x2
xsubckt_1064_nand2_x0 2 1 1535 1536 1591 nand2_x0
xsubckt_1491_nand3_x0 2 1 1163 1165 1180 1187 nand3_x0
xsubckt_153_nand2_x0 2 1 751 822 70 nand2_x0
xsubckt_170_ao22_x2 1 731 2 70 86 774 ao22_x2
xsubckt_314_a3_x2 2 570 1 691 833 20 a3_x2
xsubckt_670_nand3_x0 2 1 221 263 268 126 nand3_x0
xsubckt_719_nand3_x0 2 1 1802 263 269 138 nand3_x0
xsubckt_735_a4_x2 1 1787 2 783 831 27 20 a4_x2
xsubckt_755_a4_x2 1 1767 2 1768 1770 1771 1793 a4_x2
xsubckt_1224_oa22_x2 1 1398 2 17 528 707 oa22_x2
xsubckt_629_nand3_x0 2 1 259 263 268 129 nand3_x0
xsubckt_432_a2_x2 1 450 2 451 458 a2_x2
xsubckt_217_a2_x2 1 670 2 672 681 a2_x2
xsubckt_666_nand4_x0 2 1 224 225 226 227 228 nand4_x0
xsubckt_886_oa22_x2 1 1654 2 1657 1659 896 oa22_x2
xsubckt_1259_oa22_x2 1 1379 2 1382 1385 1393 oa22_x2
xsubckt_1497_ao22_x2 1 1157 2 1211 1170 1158 ao22_x2
xsubckt_1458_ao22_x2 1 1196 2 887 1202 1198 ao22_x2
xsubckt_482_a2_x2 1 400 2 401 402 a2_x2
xsubckt_808_oa22_x2 1 1720 2 1770 1771 850 oa22_x2
xsubckt_843_nand2_x0 2 1 1690 1769 150 nand2_x0
xsubckt_597_ao22_x2 1 290 2 715 542 484 ao22_x2
xsubckt_273_nand2_x0 2 1 611 741 747 nand2_x0
xsubckt_1039_nand4_x0 2 1 1553 784 795 20 9 nand4_x0
xsubckt_1128_nxr2_x1 1487 2 1 146 155 nxr2_x1
xsubckt_1443_a4_x2 1 1211 2 1213 1218 1222 1227 a4_x2
xsubckt_1394_nand2_x0 2 1 1257 1386 88 nand2_x0
xsubckt_1306_a3_x2 2 1336 1 1337 1346 1355 a3_x2
xsubckt_522_nand3_x0 2 1 361 570 712 800 nand3_x0
xsubckt_470_ao22_x2 1 412 2 420 416 413 ao22_x2
xsubckt_716_oa22_x2 1 185 2 288 1810 1805 oa22_x2
xsubckt_1042_a3_x2 2 1550 1 1554 741 749 a3_x2
xsubckt_1872_sff1_x4 2 202 1 1861 45 sff1_x4
xsubckt_1833_sff1_x4 2 211 1 1899 79 sff1_x4
xsubckt_1606_nand2_x0 2 1 1049 1052 1160 nand2_x0
xsubckt_1598_oa22_x2 1 1057 2 1060 1061 1188 oa22_x2
xsubckt_519_o2_x2 1 364 2 675 677 o2_x2
xsubckt_483_nand2_x0 2 1 399 401 402 nand2_x0
xsubckt_659_nand3_x0 2 1 231 263 268 127 nand3_x0
xsubckt_951_mx2_x2 1 1936 2 64 1621 553 mx2_x2
xsubckt_952_mx2_x2 1 1935 2 903 621 105 mx2_x2
xsubckt_953_mx2_x2 1 1934 2 903 628 104 mx2_x2
xsubckt_954_mx2_x2 1 1933 2 902 730 103 mx2_x2
xsubckt_1110_a2_x2 1 1902 2 1496 1505 a2_x2
xsubckt_1126_nand2_x0 2 1 1489 1490 1491 nand2_x0
xsubckt_1868_sff1_x4 2 202 1 1865 49 sff1_x4
xsubckt_1581_a3_x2 2 1074 1 1083 1085 1165 a3_x2
xsubckt_1571_a3_x2 2 1084 1 1181 1186 89 a3_x2
xsubckt_1434_a2_x2 1 1220 2 82 912 a2_x2
xsubckt_1432_oa22_x2 1 1222 2 1223 1225 883 oa22_x2
xsubckt_1404_a2_x2 1 1247 2 1248 1249 a2_x2
xsubckt_479_nand3_x0 2 1 403 405 645 767 nand3_x0
xsubckt_186_nor2_x0 2 1 708 23 20 nor2_x0
xsubckt_1060_mx2_x2 1 1538 2 747 741 761 mx2_x2
xsubckt_1209_a2_x2 1 1413 2 284 536 a2_x2
xsubckt_1829_sff1_x4 2 210 1 86 94 sff1_x4
xsubckt_1780_sff1_x4 2 208 1 1943 128 sff1_x4
xsubckt_1484_a2_x2 1 1170 2 1171 1226 a2_x2
xsubckt_136_oa22_x2 1 768 2 916 805 773 oa22_x2
xsubckt_1066_mx2_x2 1 1908 2 648 1534 81 mx2_x2
xsubckt_1776_sff1_x4 2 207 1 1947 132 sff1_x4
xsubckt_1428_oa22_x2 1 1226 2 1773 671 846 oa22_x2
xsubckt_1373_nand3_x0 2 1 1276 773 780 173 nand3_x0
xsubckt_411_nand4_x0 2 1 470 480 793 900 9 nand4_x0
xsubckt_1143_ao22_x2 1 1473 2 1474 1476 553 ao22_x2
xsubckt_1246_nand2_x0 2 1 1392 774 779 nand2_x0
xsubckt_548_nand4_x0 2 1 336 658 792 900 9 nand4_x0
xsubckt_462_nand3_x0 2 1 420 698 792 800 nand3_x0
xsubckt_60_inv_x0 2 1 165 853 inv_x0
xsubckt_243_ao22_x2 1 641 2 738 727 643 ao22_x2
xsubckt_993_nand2_x0 2 1 1592 1593 1596 nand2_x0
xsubckt_1105_nand3_x0 2 1 1500 378 619 753 nand3_x0
xsubckt_1732_oa22_x2 1 923 2 924 927 904 oa22_x2
xsubckt_1728_nxr2_x1 927 2 1 928 931 nxr2_x1
xsubckt_1574_ao22_x2 1 1081 2 1084 1086 1189 ao22_x2
xsubckt_1294_nor2_x0 2 1 1347 1348 1351 nor2_x0
xsubckt_440_oa22_x2 1 442 2 718 497 595 oa22_x2
xsubckt_61_inv_x0 2 1 164 852 inv_x0
xsubckt_62_inv_x0 2 1 163 851 inv_x0
xsubckt_63_inv_x0 2 1 162 850 inv_x0
xsubckt_64_inv_x0 2 1 161 849 inv_x0
xsubckt_65_inv_x0 2 1 67 848 inv_x0
xsubckt_66_inv_x0 2 1 65 847 inv_x0
xsubckt_174_a4_x2 1 727 2 730 747 754 760 a4_x2
xsubckt_231_nand4_x0 2 1 656 783 795 23 834 nand4_x0
xsubckt_852_nand3_x0 2 1 1683 1767 1775 54 nand3_x0
xsubckt_1746_o2_x2 1 918 2 941 904 o2_x2
xsubckt_1442_nand4_x0 2 1 1212 1214 1216 1218 1222 nand4_x0
xsubckt_621_nand4_x0 2 1 267 783 787 795 85 nand4_x0
xsubckt_67_inv_x0 2 1 35 846 inv_x0
xsubckt_68_inv_x0 2 1 94 845 inv_x0
xsubckt_69_inv_x0 2 1 192 844 inv_x0
xsubckt_192_nand3_x0 2 1 702 788 835 31 nand3_x0
xsubckt_232_a3_x2 2 655 1 656 657 663 a3_x2
xsubckt_252_a3_x2 2 632 1 681 698 719 a3_x2
xsubckt_278_nand4_x0 2 1 606 610 612 613 645 nand4_x0
xsubckt_1640_oa22_x2 1 1015 2 1160 1020 1155 oa22_x2
xsubckt_1636_nxr2_x1 1019 2 1 1031 1165 nxr2_x1
xsubckt_1366_nand2_x0 2 1 1282 1283 1289 nand2_x0
xsubckt_566_a3_x2 2 318 1 319 323 324 a3_x2
xsubckt_536_a3_x2 2 347 1 348 353 354 a3_x2
xsubckt_526_a3_x2 2 357 1 359 362 366 a3_x2
xsubckt_155_a2_x2 1 749 2 750 751 a2_x2
xsubckt_469_a2_x2 1 413 2 414 415 a2_x2
xsubckt_845_nand2_x0 2 1 1981 1689 1693 nand2_x0
xsubckt_1198_nor2_x0 2 1 1424 1425 526 nor2_x0
xsubckt_1312_ao22_x2 1 1331 2 890 1385 1333 ao22_x2
xsubckt_250_o3_x2 1 634 2 636 641 651 o3_x2
xsubckt_275_nand2_x0 2 1 609 754 760 nand2_x0
xsubckt_747_nor2_x0 2 1 1775 1776 1784 nor2_x0
xsubckt_1136_a4_x2 1 1480 2 688 719 830 886 a4_x2
xsubckt_534_o3_x2 1 349 2 350 689 797 o3_x2
xsubckt_123_o2_x2 1 790 2 16 27 o2_x2
xsubckt_1186_a4_x2 1 1436 2 784 831 27 23 a4_x2
xsubckt_1853_sff1_x4 2 207 1 1880 163 sff1_x4
xsubckt_1814_sff1_x4 2 209 1 1910 12 sff1_x4
xsubckt_1518_a3_x2 2 1137 1 1138 1139 1160 a3_x2
xsubckt_248_oa22_x2 1 636 2 692 640 637 oa22_x2
xsubckt_307_nand2_x0 2 1 577 591 794 nand2_x0
xsubckt_1888_sff1_x4 2 202 1 1845 147 sff1_x4
xsubckt_1308_mx2_x2 1 1865 2 904 1335 49 mx2_x2
xsubckt_395_nand2_x0 2 1 486 497 794 nand2_x0
xsubckt_965_nand2_x0 2 1 1930 1613 1615 nand2_x0
xsubckt_1255_ao22_x2 1 1383 2 790 565 579 ao22_x2
xsubckt_1849_sff1_x4 2 207 1 1884 167 sff1_x4
xsubckt_1761_sff1_x4 2 208 1 1956 117 sff1_x4
xsubckt_1657_mx2_x2 1 998 2 1001 1176 1189 mx2_x2
xsubckt_607_nand2_x0 2 1 281 283 633 nand2_x0
xsubckt_644_nand3_x0 2 1 245 262 268 120 nand3_x0
xsubckt_679_oa22_x2 1 188 2 288 218 1839 oa22_x2
xsubckt_1187_a2_x2 1 1435 2 479 492 a2_x2
xsubckt_1201_nand2_x0 2 1 1421 273 290 nand2_x0
xsubckt_1796_sff1_x4 2 210 1 1928 109 sff1_x4
xsubckt_1696_a2_x2 1 959 2 990 992 a2_x2
xsubckt_1647_ao22_x2 1 1008 2 241 1206 1010 ao22_x2
xsubckt_1375_nand3_x0 2 1 1274 591 793 173 nand3_x0
xsubckt_1338_nand2_x0 2 1 1308 1386 93 nand2_x0
xsubckt_554_nand3_x0 2 1 330 480 680 793 nand3_x0
xsubckt_517_nand2_x0 2 1 366 416 421 nand2_x0
xsubckt_1021_nand2_x0 2 1 1565 1566 729 nand2_x0
xsubckt_1127_xr2_x1 1488 1 2 157 156 xr2_x1
xsubckt_1268_mx2_x2 1 1869 2 903 1371 59 mx2_x2
xcmpt_mos6502_irhold_valid_hfns_2 2 1 72 69 buf_x4
xcmpt_mos6502_irhold_valid_hfns_1 2 1 69 70 buf_x4
xcmpt_mos6502_irhold_valid_hfns_0 2 1 69 71 buf_x4
xsubckt_1757_sff1_x4 2 208 1 1960 121 sff1_x4
xsubckt_1638_nand2_x0 2 1 1017 1020 1160 nand2_x0
xsubckt_1501_nand2_x0 2 1 1153 1154 1158 nand2_x0
xsubckt_1317_nxr2_x1 1326 2 1 1329 1336 nxr2_x1
xsubckt_1107_nand3_x0 2 1 1498 1499 728 755 nand3_x0
xcmpt_abc_11873_new_n561_hfns_2 2 1 649 646 buf_x4
xcmpt_abc_11873_new_n561_hfns_1 2 1 646 647 buf_x4
xcmpt_abc_11873_new_n561_hfns_0 2 1 646 648 buf_x4
xsubckt_1614_o2_x2 1 1041 2 1200 807 o2_x2
xsubckt_1555_ao22_x2 1 1100 2 1116 1118 1189 ao22_x2
xsubckt_1321_nand2_x0 2 1 1323 1325 550 nand2_x0
xsubckt_247_nand2_x0 2 1 637 638 665 nand2_x0
xsubckt_817_nand2_x0 2 1 1712 1713 1714 nand2_x0
xsubckt_1709_nxr2_x1 946 2 1 957 961 nxr2_x1
xsubckt_1444_nand4_x0 2 1 1210 1213 1218 1222 1227 nand4_x0
xsubckt_1407_nand3_x0 2 1 1245 773 780 170 nand3_x0
xsubckt_410_nand2_x0 2 1 471 480 792 nand2_x0
xsubckt_366_a4_x2 1 515 2 691 708 831 27 a4_x2
xsubckt_157_nand2_x0 2 1 744 819 70 nand2_x0
xsubckt_1264_oa22_x2 1 1374 2 153 1384 1375 oa22_x2
xsubckt_584_nand3_x0 2 1 179 302 309 433 nand3_x0
xsubckt_502_a2_x2 1 381 2 382 460 a2_x2
xsubckt_494_a3_x2 2 389 1 428 431 500 a3_x2
xsubckt_457_nand2_x0 2 1 425 515 800 nand2_x0
xsubckt_327_a2_x2 1 557 2 566 719 a2_x2
xsubckt_320_nand2_x0 2 1 564 566 832 nand2_x0
xsubckt_887_nxr2_x1 1653 2 1 1656 152 nxr2_x1
xsubckt_903_a3_x2 2 1641 1 155 160 158 a3_x2
xsubckt_923_a3_x2 2 1624 1 1663 262 268 a3_x2
xsubckt_1028_ao22_x2 1 1561 2 736 732 650 ao22_x2
xsubckt_1695_oa22_x2 1 960 2 963 966 970 oa22_x2
xsubckt_1668_nand2_x0 2 1 987 989 993 nand2_x0
xsubckt_1656_oa22_x2 1 999 2 1003 1005 1188 oa22_x2
xsubckt_1531_nand2_x0 2 1 1124 1125 1126 nand2_x0
xsubckt_562_a2_x2 1 322 2 323 324 a2_x2
xsubckt_140_nand2_x0 2 1 764 816 71 nand2_x0
xsubckt_974_nand3_x0 2 1 1606 1609 1614 621 nand3_x0
xsubckt_983_a3_x2 2 1600 1 627 731 734 a3_x2
xsubckt_1188_nand2_x0 2 1 1434 479 492 nand2_x0
xsubckt_1351_nand2_x0 2 1 1296 580 152 nand2_x0
xsubckt_620_nand2_x0 2 1 268 271 275 nand2_x0
xsubckt_706_nand3_x0 2 1 1814 263 269 139 nand3_x0
xsubckt_809_oa22_x2 1 1719 2 536 657 803 oa22_x2
xsubckt_847_nand2_x0 2 1 1687 1707 172 nand2_x0
xsubckt_1129_nxr2_x1 1486 2 1 1487 1488 nxr2_x1
xsubckt_876_a2_x2 1 1663 2 1664 9 a2_x2
xsubckt_1261_nand2_x0 2 1 1377 1380 579 nand2_x0
xcmpt_mos6502_state_bit4_hfns_2 2 1 28 15 buf_x4
xcmpt_mos6502_state_bit4_hfns_1 2 1 15 16 buf_x4
xcmpt_mos6502_state_bit4_hfns_0 2 1 15 17 buf_x4
xcmpt_mos6502_state_bit3_hfns_2 2 1 29 18 buf_x4
xcmpt_mos6502_state_bit3_hfns_1 2 1 18 19 buf_x4
xcmpt_mos6502_state_bit3_hfns_0 2 1 18 20 buf_x4
xcmpt_mos6502_state_bit2_hfns_2 2 1 30 21 buf_x4
xcmpt_mos6502_state_bit2_hfns_1 2 1 21 22 buf_x4
xcmpt_mos6502_state_bit2_hfns_0 2 1 21 23 buf_x4
xcmpt_mos6502_state_bit0_hfns_2 2 1 32 24 buf_x4
xcmpt_mos6502_state_bit0_hfns_1 2 1 24 25 buf_x4
xcmpt_mos6502_state_bit0_hfns_0 2 1 24 26 buf_x4
xsubckt_1873_sff1_x4 2 206 1 1860 44 sff1_x4
xsubckt_1724_ao22_x2 1 931 2 933 934 1119 ao22_x2
xsubckt_1398_a4_x2 1 1253 2 1254 1255 1256 549 a4_x2
xsubckt_260_nand2_x0 2 1 624 837 71 nand2_x0
xsubckt_804_o2_x2 1 1973 2 1724 1731 o2_x2
xsubckt_830_nand2_x0 2 1 1701 1780 92 nand2_x0
xsubckt_960_mx2_x2 1 1616 2 647 627 43 mx2_x2
xsubckt_1834_sff1_x4 2 211 1 1898 78 sff1_x4
xsubckt_1671_a3_x2 2 984 1 1181 1186 93 a3_x2
xsubckt_1651_a3_x2 2 1004 1 1181 1186 92 a3_x2
xsubckt_1420_nand3_x0 2 1 1233 591 794 169 nand3_x0
xsubckt_346_nand3_x0 2 1 535 543 713 800 nand3_x0
xsubckt_664_oa22_x2 1 226 2 253 700 893 oa22_x2
xsubckt_874_o2_x2 1 1665 2 1787 668 o2_x2
xsubckt_1012_o4_x2 1 1573 2 1576 1582 1588 1592 o4_x2
xsubckt_1055_a2_x2 1 1541 2 1600 621 a2_x2
xsubckt_1075_a2_x2 1 1525 2 1526 650 a2_x2
xsubckt_1115_mx2_x2 1 1900 2 1495 93 80 mx2_x2
xsubckt_1116_mx2_x2 1 1899 2 1495 92 79 mx2_x2
xsubckt_1260_a2_x2 1 1378 2 1380 579 a2_x2
xsubckt_1869_sff1_x4 2 202 1 1864 48 sff1_x4
xsubckt_1781_sff1_x4 2 208 1 1942 127 sff1_x4
xsubckt_1564_a2_x2 1 1091 2 1102 1227 a2_x2
xsubckt_1557_nand3_x0 2 1 1098 1115 1117 1176 nand3_x0
xsubckt_1544_a2_x2 1 1111 2 1113 1160 a2_x2
xsubckt_1524_a2_x2 1 1131 2 1132 1133 a2_x2
xsubckt_1467_nand3_x0 2 1 1187 698 793 46 nand3_x0
xsubckt_176_oa22_x2 1 725 2 726 737 767 oa22_x2
xsubckt_1085_a2_x2 1 1906 2 1517 1523 a2_x2
xsubckt_1117_mx2_x2 1 1898 2 1495 91 78 mx2_x2
xsubckt_1118_mx2_x2 1 1897 2 1495 90 77 mx2_x2
xsubckt_1119_mx2_x2 1 1896 2 1495 89 76 mx2_x2
xsubckt_1429_oa22_x2 1 1225 2 1773 671 879 oa22_x2
xsubckt_1399_a2_x2 1 1252 2 1253 1257 a2_x2
xsubckt_1389_a2_x2 1 1261 2 1262 1267 a2_x2
xsubckt_646_nand3_x0 2 1 243 263 269 144 nand3_x0
xsubckt_1113_nand2_x0 2 1 1493 1494 648 nand2_x0
xsubckt_1150_nand3_x0 2 1 1468 585 700 777 nand3_x0
xsubckt_1777_sff1_x4 2 208 1 1946 131 sff1_x4
xsubckt_1540_nand3_x0 2 1 1115 1181 1186 88 nand3_x0
xsubckt_593_nand4_x0 2 1 293 591 680 831 27 nand4_x0
xsubckt_860_nand2_x0 2 1 1676 1780 87 nand2_x0
xsubckt_1413_nand2_x0 2 1 1239 1241 1246 nand2_x0
xsubckt_529_oa22_x2 1 354 2 371 372 644 oa22_x2
xsubckt_70_inv_x0 2 1 73 843 inv_x0
xsubckt_71_inv_x0 2 1 95 842 inv_x0
xsubckt_72_inv_x0 2 1 193 841 inv_x0
xsubckt_73_inv_x0 2 1 74 840 inv_x0
xsubckt_205_ao22_x2 1 686 2 710 687 689 ao22_x2
xsubckt_715_nand4_x0 2 1 1805 1806 1807 1808 1809 nand4_x0
xsubckt_819_nand2_x0 2 1 1710 1711 1716 nand2_x0
xsubckt_1729_nxr2_x1 926 2 1 935 937 nxr2_x1
xsubckt_1409_nand3_x0 2 1 1243 591 792 170 nand3_x0
xsubckt_1319_nand3_x0 2 1 1325 773 780 162 nand3_x0
xsubckt_568_a4_x2 1 316 2 317 410 465 598 a4_x2
xsubckt_558_a4_x2 1 326 2 327 394 403 406 a4_x2
xsubckt_74_inv_x0 2 1 96 839 inv_x0
xsubckt_75_inv_x0 2 1 194 838 inv_x0
xsubckt_76_inv_x0 2 1 75 837 inv_x0
xsubckt_77_inv_x0 2 1 31 836 inv_x0
xsubckt_78_inv_x0 2 1 26 835 inv_x0
xsubckt_79_inv_x0 2 1 20 834 inv_x0
xsubckt_1270_nand3_x0 2 1 1369 773 780 167 nand3_x0
xsubckt_578_a4_x2 1 307 2 561 567 602 603 a4_x2
xsubckt_322_nand2_x0 2 1 562 566 713 nand2_x0
xsubckt_177_a3_x2 2 724 1 788 26 836 a3_x2
xsubckt_187_a3_x2 2 707 1 708 26 836 a3_x2
xsubckt_225_a2_x2 1 662 2 17 27 a2_x2
xsubckt_811_a3_x2 2 1717 1 1718 1721 1722 a3_x2
xsubckt_1002_nand3_x0 2 1 1583 1585 1587 753 nand3_x0
xsubckt_1053_nand2_x0 2 1 1542 1543 1544 nand2_x0
xsubckt_1676_oa22_x2 1 979 2 1160 981 1155 oa22_x2
xsubckt_1570_nand3_x0 2 1 1085 698 795 49 nand3_x0
xsubckt_460_a2_x2 1 422 2 423 427 a2_x2
xsubckt_369_nand2_x0 2 1 512 515 681 nand2_x0
xsubckt_148_ao22_x2 1 756 2 71 90 774 ao22_x2
xsubckt_265_a2_x2 1 619 2 729 766 a2_x2
xsubckt_1480_nand3_x0 2 1 1174 1177 1190 1192 nand3_x0
xsubckt_579_a2_x2 1 306 2 307 308 a2_x2
xsubckt_549_a2_x2 1 335 2 336 337 a2_x2
xsubckt_702_oa22_x2 1 1817 2 486 568 873 oa22_x2
xsubckt_708_nand3_x0 2 1 1812 263 268 123 nand3_x0
xsubckt_744_a2_x2 1 1778 2 530 539 a2_x2
xsubckt_849_nand2_x0 2 1 1685 1769 149 nand2_x0
xsubckt_1421_a4_x2 1 1232 2 1233 1234 1235 549 a4_x2
xsubckt_390_o3_x2 1 491 2 492 797 832 o3_x2
xsubckt_175_nand4_x0 2 1 726 730 747 754 760 nand4_x0
xsubckt_213_o2_x2 1 674 2 675 797 o2_x2
xsubckt_1030_a3_x2 2 1559 1 729 742 747 a3_x2
xsubckt_1702_mx2_x2 1 953 2 1021 1016 1018 mx2_x2
xsubckt_1296_a4_x2 1 1345 2 1346 1356 1364 1373 a4_x2
xsubckt_537_o2_x2 1 346 2 539 797 o2_x2
xsubckt_211_nand3_x0 2 1 676 681 722 27 nand3_x0
xsubckt_1090_a3_x2 2 1512 1 1513 1514 1583 a3_x2
xsubckt_1854_sff1_x4 2 202 1 1879 162 sff1_x4
xsubckt_1815_sff1_x4 2 205 1 1909 14 sff1_x4
xsubckt_1563_nand2_x0 2 1 1092 1094 1108 nand2_x0
xsubckt_1492_oa22_x2 1 1162 2 1187 1180 1165 oa22_x2
xsubckt_1412_a2_x2 1 1240 2 1241 1246 a2_x2
xsubckt_601_nand3_x0 2 1 286 655 694 705 nand3_x0
xsubckt_475_nand4_x0 2 1 407 610 645 740 767 nand4_x0
xsubckt_385_nand4_x0 2 1 496 833 20 26 836 nand4_x0
xsubckt_172_nand2_x0 2 1 729 733 735 nand2_x0
xsubckt_262_nand2_x0 2 1 622 624 774 nand2_x0
xsubckt_828_nand3_x0 2 1 1703 1767 1775 44 nand3_x0
xsubckt_969_nand2_x0 2 1 1610 648 109 nand2_x0
xsubckt_1079_nand3_x0 2 1 1522 1575 378 609 nand3_x0
xsubckt_1199_a3_x2 2 1423 1 1424 1426 1428 a3_x2
xsubckt_1889_sff1_x4 2 202 1 1844 146 sff1_x4
xsubckt_1762_sff1_x4 2 207 1 1955 116 sff1_x4
xsubckt_1706_a2_x2 1 949 2 672 160 a2_x2
xsubckt_1663_mx2_x2 1 992 2 1227 995 1037 mx2_x2
xsubckt_1662_mx2_x2 1 993 2 1227 994 1036 mx2_x2
xsubckt_1661_mx2_x2 1 994 2 1008 996 1000 mx2_x2
xsubckt_1660_mx2_x2 1 995 2 1008 997 999 mx2_x2
xsubckt_1613_ao22_x2 1 1042 2 1203 1789 151 ao22_x2
xsubckt_1482_a2_x2 1 1172 2 1173 1174 a2_x2
xsubckt_1472_a2_x2 1 1182 2 1407 1438 a2_x2
xsubckt_1452_a2_x2 1 1202 2 1204 1790 a2_x2
xsubckt_1383_nand2_x0 2 1 1267 1379 55 nand2_x0
xsubckt_1318_mx2_x2 1 1864 2 903 1326 48 mx2_x2
xsubckt_129_nor2_x0 2 1 775 177 64 nor2_x0
xsubckt_738_nand3_x0 2 1 1784 1786 1788 1790 nand3_x0
xsubckt_1687_ao22_x2 1 968 2 1167 1166 1161 ao22_x2
xsubckt_599_nor2_x0 2 1 288 289 701 nor2_x0
xsubckt_685_nand4_x0 2 1 1833 1835 1836 1837 1838 nand4_x0
xsubckt_1277_mx2_x2 1 1868 2 904 1363 58 mx2_x2
xsubckt_417_nand4_x0 2 1 464 466 498 509 516 nand4_x0
xsubckt_468_nand3_x0 2 1 414 591 680 831 nand3_x0
xsubckt_1357_nxr2_x1 1290 2 1 1292 1300 nxr2_x1
xsubckt_1797_sff1_x4 2 210 1 1927 38 sff1_x4
xsubckt_1758_sff1_x4 2 208 1 1959 120 sff1_x4
xsubckt_999_nand2_x0 2 1 1586 1587 753 nand2_x0
xsubckt_858_nand3_x0 2 1 1678 1767 1775 53 nand3_x0
xsubckt_416_a4_x2 1 465 2 466 498 509 516 a4_x2
xsubckt_611_a4_x2 1 277 2 521 553 667 675 a4_x2
xsubckt_1295_o2_x2 1 1346 2 1348 1351 o2_x2
xsubckt_1679_nand3_x0 2 1 976 983 985 1176 nand3_x0
xsubckt_892_nxr2_x1 1649 2 1 1660 893 nxr2_x1
xsubckt_288_nand3_x0 2 1 596 691 23 834 nand3_x0
xsubckt_504_nand2_x0 2 1 379 380 437 nand2_x0
xsubckt_1362_nand3_x0 2 1 1286 591 795 174 nand3_x0
xsubckt_982_nand2_x0 2 1 1601 648 107 nand2_x0
xsubckt_143_a2_x2 1 761 2 763 765 a2_x2
xsubckt_359_a3_x2 2 522 1 658 17 832 a3_x2
xsubckt_451_nand3_x0 2 1 431 462 612 753 nand3_x0
xsubckt_514_a3_x2 2 369 1 370 404 435 a3_x2
xsubckt_1625_nand2_x0 2 1 1030 1032 1034 nand2_x0
xsubckt_838_a3_x2 2 1694 1 1695 1696 1697 a3_x2
xsubckt_220_nand4_x0 2 1 667 784 788 17 832 nand4_x0
xsubckt_193_a2_x2 1 701 2 703 719 a2_x2
xsubckt_183_a2_x2 1 714 2 17 832 a2_x2
xsubckt_144_nand2_x0 2 1 760 763 765 nand2_x0
xsubckt_437_a2_x2 1 445 2 688 719 a2_x2
xsubckt_594_a3_x2 2 292 1 293 294 331 a3_x2
xsubckt_1572_nand3_x0 2 1 1083 1181 1186 89 nand3_x0
xsubckt_868_a3_x2 2 1669 1 1670 1671 1672 a3_x2
xsubckt_520_nand4_x0 2 1 363 681 784 788 794 nand4_x0
xsubckt_1124_nand3_x0 2 1 1491 1492 585 777 nand3_x0
xsubckt_206_nor2_x0 2 1 685 14 155 nor2_x0
xsubckt_430_nand4_x0 2 1 452 454 610 612 645 nand4_x0
xsubckt_1745_nand2_x0 2 1 919 154 904 nand2_x0
xsubckt_956_ao22_x2 1 1619 2 773 630 650 ao22_x2
xsubckt_340_nand4_x0 2 1 541 708 794 835 31 nand4_x0
xsubckt_481_nand3_x0 2 1 401 566 679 794 nand3_x0
xsubckt_625_mx2_x2 1 263 2 270 265 829 mx2_x2
xsubckt_1468_a4_x2 1 1186 2 1404 1418 519 583 a4_x2
xsubckt_1800_sff1_x4 2 210 1 1924 107 sff1_x4
xsubckt_1122_mx2_x2 1 1893 2 1495 86 73 mx2_x2
xsubckt_1121_mx2_x2 1 1894 2 1495 87 74 mx2_x2
xsubckt_1120_mx2_x2 1 1895 2 1495 88 75 mx2_x2
xsubckt_957_nand4_x0 2 1 1618 1619 462 612 753 nand4_x0
xsubckt_665_oa22_x2 1 225 2 249 550 917 oa22_x2
xsubckt_650_o2_x2 1 239 2 256 864 o2_x2
xsubckt_264_nand2_x0 2 1 620 623 625 nand2_x0
xsubckt_626_mx2_x2 1 262 2 270 264 34 mx2_x2
xsubckt_1300_a2_x2 1 1342 2 1343 550 a2_x2
xsubckt_1310_a2_x2 1 1333 2 1334 550 a2_x2
xsubckt_1320_a2_x2 1 1324 2 1325 550 a2_x2
xsubckt_1565_nand2_x0 2 1 1090 1102 1227 nand2_x0
xsubckt_1835_sff1_x4 2 211 1 1897 77 sff1_x4
xsubckt_1874_sff1_x4 2 206 1 1859 57 sff1_x4
xsubckt_1195_a2_x2 1 1427 2 589 700 a2_x2
xsubckt_825_ao22_x2 1 1705 2 897 1770 1793 ao22_x2
xsubckt_1370_a2_x2 1 1278 2 1279 1280 a2_x2
xsubckt_1381_nxr2_x1 1268 2 1 1271 1281 nxr2_x1
xsubckt_1475_nand2_x0 2 1 1179 1180 1187 nand2_x0
xsubckt_1624_a2_x2 1 1031 2 1032 1034 a2_x2
xsubckt_1184_ao22_x2 1 1438 2 715 687 667 ao22_x2
xsubckt_423_nand3_x0 2 1 459 461 610 612 nand3_x0
xsubckt_1469_a2_x2 1 1185 2 290 507 a2_x2
xsubckt_1782_sff1_x4 2 208 1 1941 126 sff1_x4
xsubckt_1106_ao22_x2 1 1499 2 622 626 627 ao22_x2
xsubckt_1027_nand2_x0 2 1 1562 648 40 nand2_x0
xsubckt_1013_nand4_x0 2 1 1572 455 729 741 749 nand4_x0
xsubckt_813_nand3_x0 2 1 1716 1767 1775 46 nand3_x0
xsubckt_1303_oa22_x2 1 1339 2 149 1384 1341 oa22_x2
xsubckt_1507_nand2_x0 2 1 1148 1149 1306 nand2_x0
xsubckt_1778_sff1_x4 2 206 1 1945 130 sff1_x4
xsubckt_304_a4_x2 1 580 2 691 792 23 834 a4_x2
xsubckt_80_inv_x0 2 1 22 833 inv_x0
xsubckt_1417_nand2_x0 2 1 1236 1379 52 nand2_x0
xsubckt_1447_o2_x2 1 1207 2 1209 1224 o2_x2
xsubckt_1502_ao22_x2 1 1152 2 1155 1159 9 ao22_x2
xsubckt_1584_o3_x2 1 1071 2 1073 1074 1161 o3_x2
xsubckt_1100_nand2_x0 2 1 1505 647 848 nand2_x0
xsubckt_179_a4_x2 1 722 2 787 831 26 836 a4_x2
xsubckt_81_inv_x0 2 1 27 832 inv_x0
xsubckt_82_inv_x0 2 1 17 831 inv_x0
xsubckt_83_inv_x0 2 1 37 830 inv_x0
xsubckt_84_inv_x0 2 1 34 829 inv_x0
xsubckt_85_inv_x0 2 1 85 828 inv_x0
xsubckt_86_inv_x0 2 1 81 827 inv_x0
xsubckt_384_a4_x2 1 497 2 833 20 25 836 a4_x2
xsubckt_618_a4_x2 1 270 2 272 276 282 777 a4_x2
xsubckt_1734_oa22_x2 1 922 2 969 963 966 oa22_x2
xsubckt_1133_nand4_x0 2 1 1482 1483 784 788 795 nand4_x0
xsubckt_1006_nand3_x0 2 1 1579 1609 620 766 nand3_x0
xsubckt_698_a4_x2 1 1821 2 1823 1824 1825 1826 a4_x2
xsubckt_648_a4_x2 1 241 2 242 243 244 245 a4_x2
xsubckt_287_a3_x2 2 597 1 691 23 834 a3_x2
xsubckt_277_a3_x2 2 607 1 610 612 613 a3_x2
xsubckt_267_a3_x2 2 617 1 620 729 766 a3_x2
xsubckt_87_inv_x0 2 1 33 826 inv_x0
xsubckt_88_inv_x0 2 1 84 825 inv_x0
xsubckt_89_inv_x0 2 1 101 824 inv_x0
xsubckt_363_nand3_x0 2 1 518 528 800 17 nand3_x0
xsubckt_472_a3_x2 2 410 1 411 433 450 a3_x2
xsubckt_500_a2_x2 1 383 2 384 725 a2_x2
xsubckt_1400_nand2_x0 2 1 1251 1252 1258 nand2_x0
xsubckt_1603_nxr2_x1 1052 2 1 1059 1164 nxr2_x1
xsubckt_941_a3_x2 2 1622 1 1663 263 268 a3_x2
xsubckt_753_nand3_x0 2 1 1769 579 656 694 nand3_x0
xsubckt_736_a3_x2 2 1786 1 521 568 585 a3_x2
xsubckt_550_a2_x2 1 334 2 335 338 a2_x2
xsubckt_609_a2_x2 1 279 2 521 553 a2_x2
xsubckt_637_ao22_x2 1 251 2 543 703 719 ao22_x2
xsubckt_1688_nor2_x0 2 1 967 968 1227 nor2_x0
xsubckt_146_nand2_x0 2 1 758 813 71 nand2_x0
xsubckt_570_a2_x2 1 314 2 315 545 a2_x2
xsubckt_619_a2_x2 1 269 2 271 275 a2_x2
xsubckt_1040_nand2_x0 2 1 1552 1553 160 nand2_x0
xsubckt_884_a2_x2 1 1656 2 1657 1659 a2_x2
xsubckt_1314_ao22_x2 1 1329 2 873 1378 1331 ao22_x2
xsubckt_1316_a4_x2 1 1327 2 1328 1337 1346 1355 a4_x2
xsubckt_1747_nand2_x0 2 1 1843 918 919 nand2_x0
xsubckt_1036_nand3_x0 2 1 1555 1556 1577 650 nand3_x0
xsubckt_912_nand4_x0 2 1 1633 147 155 160 158 nand4_x0
xsubckt_836_nand2_x0 2 1 1696 1769 151 nand2_x0
xsubckt_802_o2_x2 1 1725 2 1726 1729 o2_x2
xsubckt_128_o2_x2 1 776 2 89 71 o2_x2
xsubckt_342_nand4_x0 2 1 539 691 708 17 832 nand4_x0
xsubckt_343_o2_x2 1 538 2 539 677 o2_x2
xsubckt_393_nand3_x0 2 1 488 494 713 800 nand3_x0
xsubckt_1346_a4_x2 1 1300 2 1301 1314 1319 1327 a4_x2
xsubckt_1376_a4_x2 1 1273 2 1274 1275 1276 549 a4_x2
xsubckt_1388_ao22_x2 1 1262 2 805 1387 1263 ao22_x2
xsubckt_1820_sff1_x4 2 209 1 1904 84 sff1_x4
xsubckt_1249_a3_x2 2 1389 1 1390 502 541 a3_x2
xsubckt_1087_nand2_x0 2 1 1515 760 767 nand2_x0
xsubckt_1063_a2_x2 1 1536 2 1600 767 a2_x2
xsubckt_266_nand2_x0 2 1 618 729 766 nand2_x0
xsubckt_389_nand4_x0 2 1 492 784 831 833 20 nand4_x0
xsubckt_605_nand3_x0 2 1 283 566 661 790 nand3_x0
xsubckt_1415_nxr2_x1 1237 2 1 1240 1250 nxr2_x1
xsubckt_1439_nor3_x0 2 1 1215 1410 537 557 nor3_x0
xsubckt_1516_nand3_x0 2 1 1139 1140 1142 1165 nand3_x0
xsubckt_1816_sff1_x4 2 209 1 1908 81 sff1_x4
xsubckt_1855_sff1_x4 2 206 1 1878 161 sff1_x4
xsubckt_1218_ao22_x2 1 1404 2 715 596 530 ao22_x2
xsubckt_1109_o4_x2 1 1496 2 1497 1501 1503 1519 o4_x2
xsubckt_1093_a2_x2 1 1510 2 648 825 a2_x2
xsubckt_1058_oa22_x2 1 1910 2 1599 1544 1540 oa22_x2
xsubckt_693_nand3_x0 2 1 1826 263 268 124 nand3_x0
xsubckt_642_nand4_x0 2 1 246 247 250 254 255 nand4_x0
xsubckt_1327_mx2_x2 1 1863 2 903 1318 47 mx2_x2
xsubckt_1532_a2_x2 1 1123 2 1124 1174 a2_x2
xsubckt_425_nand3_x0 2 1 457 566 680 718 nand3_x0
xsubckt_1550_nand2_x0 2 1 1105 1107 1255 nand2_x0
xsubckt_1763_sff1_x4 2 207 1 1954 115 sff1_x4
xsubckt_1015_nand4_x0 2 1 1570 620 729 741 749 nand4_x0
xsubckt_866_nand2_x0 2 1 1671 1780 86 nand2_x0
xsubckt_245_nand3_x0 2 1 639 685 900 9 nand3_x0
xsubckt_1289_mx2_x2 1 1867 2 904 1352 51 mx2_x2
xsubckt_1323_oa22_x2 1 1321 2 147 1384 1323 oa22_x2
xsubckt_1798_sff1_x4 2 210 1 1926 108 sff1_x4
xsubckt_282_nand4_x0 2 1 602 684 688 712 800 nand4_x0
xsubckt_222_a4_x2 1 665 2 666 669 674 676 a4_x2
xsubckt_635_nand3_x0 2 1 253 543 719 866 nand3_x0
xsubckt_1419_nand2_x0 2 1 1234 580 146 nand2_x0
xsubckt_1597_nand2_x0 2 1 1058 1060 1061 nand2_x0
xsubckt_1759_sff1_x4 2 210 1 1958 119 sff1_x4
xsubckt_1280_nand2_x0 2 1 1360 64 915 nand2_x0
xsubckt_1190_nand2_x0 2 1 1432 541 667 nand2_x0
xsubckt_893_nxr2_x1 1648 2 1 1649 1654 nxr2_x1
xsubckt_749_ao22_x2 1 1773 2 715 687 514 ao22_x2
xsubckt_741_a4_x2 1 1781 2 1783 593 664 686 a4_x2
xsubckt_721_a4_x2 1 1800 2 1801 1802 1803 1804 a4_x2
xsubckt_310_a3_x2 2 574 1 576 900 9 a3_x2
xsubckt_404_nand4_x0 2 1 477 480 662 900 9 nand4_x0
xsubckt_508_nand2_x0 2 1 375 376 377 nand2_x0
xsubckt_545_nand3_x0 2 1 339 480 662 681 nand3_x0
xsubckt_622_ao22_x2 1 266 2 827 272 267 ao22_x2
xsubckt_1329_nand2_x0 2 1 1316 1317 550 nand2_x0
xsubckt_1609_o2_x2 1 1046 2 1048 1053 o2_x2
xsubckt_1008_nand3_x0 2 1 1577 1581 612 752 nand3_x0
xsubckt_986_nand2_x0 2 1 1924 1598 1601 nand2_x0
xsubckt_586_a4_x2 1 300 2 452 457 503 506 a4_x2
xsubckt_1580_nand2_x0 2 1 1075 1077 1080 nand2_x0
xsubckt_1227_oa22_x2 1 1395 2 1396 1422 903 oa22_x2
xsubckt_1059_nand2_x0 2 1 1539 648 14 nand2_x0
xsubckt_815_oa22_x2 1 1714 2 536 657 802 oa22_x2
xsubckt_263_a2_x2 1 621 2 623 625 a2_x2
xsubckt_224_nand4_x0 2 1 663 708 795 26 836 nand4_x0
xsubckt_449_a3_x2 2 433 1 434 439 440 a3_x2
xsubckt_459_a3_x2 2 423 1 424 425 426 a3_x2
xsubckt_507_a2_x2 1 376 2 438 766 a2_x2
xsubckt_614_nand4_x0 2 1 274 784 788 794 84 nand4_x0
xsubckt_998_a3_x2 2 1587 1 741 747 766 a3_x2
xsubckt_961_ao22_x2 1 1931 2 647 505 1616 ao22_x2
xsubckt_723_oa22_x2 1 1798 2 486 568 871 oa22_x2
xsubckt_221_nand2_x0 2 1 666 668 800 nand2_x0
xsubckt_580_nor4_x0 2 1 305 358 472 487 587 nor4_x0
xsubckt_1359_nand2_x0 2 1 1289 1379 57 nand2_x0
xsubckt_1396_nand3_x0 2 1 1255 591 794 171 nand3_x0
xsubckt_1619_oa22_x2 1 1036 2 229 1205 1038 oa22_x2
xsubckt_758_oa22_x2 1 1764 2 1770 1771 856 oa22_x2
xsubckt_701_nand2_x0 2 1 1818 251 148 nand2_x0
xsubckt_700_o2_x2 1 1819 2 256 859 o2_x2
xsubckt_235_oa22_x2 1 652 2 655 659 797 oa22_x2
xsubckt_485_nand3_x0 2 1 397 543 680 718 nand3_x0
xsubckt_1332_a3_x2 2 1313 1 1314 1319 1327 a3_x2
xsubckt_1659_nand2_x0 2 1 996 998 1174 nand2_x0
xsubckt_1801_sff1_x4 2 209 1 1923 112 sff1_x4
xsubckt_1840_sff1_x4 2 210 1 1892 13 sff1_x4
xsubckt_918_ao22_x2 1 1628 2 1636 1632 1633 ao22_x2
xsubckt_734_nand4_x0 2 1 1788 783 831 27 20 nand4_x0
xsubckt_127_nand3_x0 2 1 777 783 788 793 nand3_x0
xsubckt_575_o2_x2 1 180 2 310 316 o2_x2
xsubckt_1527_oa22_x2 1 1128 2 1810 1205 1130 oa22_x2
xsubckt_1875_sff1_x4 2 206 1 1858 56 sff1_x4
xsubckt_1245_a2_x2 1 1393 2 774 779 a2_x2
xsubckt_1135_mx2_x2 1 1892 2 1489 1481 13 mx2_x2
xsubckt_695_nand3_x0 2 1 1824 263 269 140 nand3_x0
xsubckt_164_nand4_x0 2 1 737 741 749 755 760 nand4_x0
xsubckt_1430_a2_x2 1 1224 2 672 880 a2_x2
xsubckt_1440_a2_x2 1 1214 2 1215 1217 a2_x2
xsubckt_1836_sff1_x4 2 209 1 1896 76 sff1_x4
xsubckt_1138_mx2_x2 1 1478 2 780 585 909 mx2_x2
xsubckt_989_mx2_x2 1 1923 2 648 1597 112 mx2_x2
xsubckt_251_nand2_x0 2 1 633 697 719 nand2_x0
xsubckt_427_nand3_x0 2 1 455 623 625 628 nand3_x0
xsubckt_478_nand2_x0 2 1 404 405 767 nand2_x0
xsubckt_585_nor2_x0 2 1 301 510 604 nor2_x0
xsubckt_1481_mx2_x2 1 1173 2 1179 1176 1189 mx2_x2
xsubckt_1483_mx2_x2 1 1171 2 1194 1172 1178 mx2_x2
xsubckt_1559_a2_x2 1 1096 2 1097 1174 a2_x2
xsubckt_1579_a2_x2 1 1076 2 1077 1080 a2_x2
xsubckt_1783_sff1_x4 2 207 1 1940 125 sff1_x4
xsubckt_958_nand2_x0 2 1 1932 1618 1620 nand2_x0
xsubckt_778_nand2_x0 2 1 1746 1747 1752 nand2_x0
xsubckt_219_a4_x2 1 668 2 784 788 16 832 a4_x2
xsubckt_1372_nand2_x0 2 1 1277 1379 56 nand2_x0
xsubckt_1700_oa22_x2 1 955 2 958 960 988 oa22_x2
xsubckt_1779_sff1_x4 2 208 1 1944 129 sff1_x4
xsubckt_1104_nand2_x0 2 1 1501 1502 1586 nand2_x0
xsubckt_229_a4_x2 1 658 2 23 20 26 31 a4_x2
xsubckt_90_inv_x0 2 1 199 823 inv_x0
xsubckt_91_inv_x0 2 1 80 822 inv_x0
xsubckt_92_inv_x0 2 1 100 821 inv_x0
xsubckt_93_inv_x0 2 1 198 820 inv_x0
xsubckt_444_a4_x2 1 438 2 756 758 762 764 a4_x2
xsubckt_1368_nand3_x0 2 1 1280 1282 1291 1300 nand3_x0
xsubckt_1621_nand3_x0 2 1 1034 698 795 51 nand3_x0
xsubckt_1170_nor2_x0 2 1 1450 42 110 nor2_x0
xsubckt_1137_nand4_x0 2 1 1479 688 719 830 886 nand4_x0
xsubckt_851_nand2_x0 2 1 1980 1684 1688 nand2_x0
xsubckt_800_oa22_x2 1 1727 2 1770 1771 851 oa22_x2
xsubckt_289_a4_x2 1 595 2 691 832 23 834 a4_x2
xsubckt_230_nand3_x0 2 1 657 658 831 27 nand3_x0
xsubckt_94_inv_x0 2 1 79 819 inv_x0
xsubckt_95_inv_x0 2 1 99 818 inv_x0
xsubckt_96_inv_x0 2 1 197 817 inv_x0
xsubckt_97_inv_x0 2 1 78 816 inv_x0
xsubckt_98_inv_x0 2 1 98 815 inv_x0
xsubckt_99_inv_x0 2 1 196 814 inv_x0
xsubckt_141_a2_x2 1 763 2 764 774 a2_x2
xsubckt_1411_ao22_x2 1 1241 2 803 1387 1242 ao22_x2
xsubckt_1587_o2_x2 1 1068 2 1200 806 o2_x2
xsubckt_963_a4_x2 1 1614 2 612 650 753 767 a4_x2
xsubckt_181_a2_x2 1 720 2 831 27 a2_x2
xsubckt_171_a2_x2 1 730 2 733 735 a2_x2
xsubckt_161_a2_x2 1 740 2 741 749 a2_x2
xsubckt_151_a2_x2 1 753 2 755 760 a2_x2
xsubckt_154_ao22_x2 1 750 2 71 93 774 ao22_x2
xsubckt_387_a3_x2 2 494 1 784 833 20 a3_x2
xsubckt_402_o4_x2 1 479 2 23 20 26 31 o4_x2
xsubckt_572_a3_x2 2 312 1 451 458 516 a3_x2
xsubckt_1604_nxr2_x1 1051 2 1 1059 1165 nxr2_x1
xsubckt_1682_oa22_x2 1 973 2 976 977 1175 oa22_x2
xsubckt_856_a3_x2 2 1679 1 1680 1681 1682 a3_x2
xsubckt_403_nand2_x0 2 1 478 480 662 nand2_x0
xsubckt_530_nand3_x0 2 1 353 679 688 718 nand3_x0
xsubckt_640_a2_x2 1 248 2 249 550 a2_x2
xsubckt_1155_oa22_x2 1 1463 2 703 718 780 oa22_x2
xsubckt_782_oa22_x2 1 1743 2 1770 1771 853 oa22_x2
xsubckt_769_a2_x2 1 1754 2 1755 1756 a2_x2
xsubckt_704_oa22_x2 1 186 2 288 1820 1816 oa22_x2
xsubckt_546_ao22_x2 1 338 2 532 393 339 ao22_x2
xsubckt_1354_ao22_x2 1 1293 2 808 1387 1294 ao22_x2
xsubckt_1678_oa22_x2 1 977 2 983 985 1188 oa22_x2
xsubckt_1200_a3_x2 2 1422 1 1423 1430 1433 a3_x2
xsubckt_1005_a3_x2 2 1580 1 1609 620 766 a3_x2
xsubckt_967_nand3_x0 2 1 1611 1614 355 621 nand3_x0
xsubckt_133_nand2_x0 2 1 771 810 71 nand2_x0
xsubckt_1821_sff1_x4 2 205 1 1903 41 sff1_x4
xsubckt_1860_sff1_x4 2 206 1 1873 172 sff1_x4
xsubckt_1262_ao22_x2 1 1376 2 1379 580 59 ao22_x2
xsubckt_1223_ao22_x2 1 1399 2 1422 1411 1400 ao22_x2
xsubckt_739_oa22_x2 1 1783 2 715 710 496 oa22_x2
xsubckt_651_oa22_x2 1 238 2 486 568 877 oa22_x2
xsubckt_523_nand2_x0 2 1 360 668 680 nand2_x0
xsubckt_1514_a3_x2 2 1141 1 1181 1186 87 a3_x2
xsubckt_1547_oa22_x2 1 1108 2 1160 1113 1155 oa22_x2
xsubckt_1720_mx2_x2 1 935 2 1093 1109 1111 mx2_x2
xsubckt_697_nand3_x0 2 1 1822 1823 1824 1825 nand3_x0
xsubckt_308_xr2_x1 576 1 2 113 155 xr2_x1
xsubckt_560_nand3_x0 2 1 324 494 680 712 nand3_x0
xsubckt_1291_nand3_x0 2 1 1350 773 780 165 nand3_x0
xsubckt_1336_mx2_x2 1 1862 2 904 1310 46 mx2_x2
xsubckt_1494_oa22_x2 1 1160 2 1773 671 867 oa22_x2
xsubckt_1723_mx2_x2 1 932 2 1120 1135 1137 mx2_x2
xsubckt_1817_sff1_x4 2 210 1 1907 34 sff1_x4
xsubckt_1856_sff1_x4 2 202 1 1877 176 sff1_x4
xsubckt_1258_ao22_x2 1 1380 2 1381 1384 1392 ao22_x2
xsubckt_885_ao22_x2 1 1655 2 1658 1660 152 ao22_x2
xsubckt_202_nand3_x0 2 1 689 691 708 792 nand3_x0
xsubckt_380_nand3_x0 2 1 501 680 697 792 nand3_x0
xsubckt_429_nand3_x0 2 1 453 456 729 766 nand3_x0
xsubckt_1644_nand2_x0 2 1 1011 1012 1295 nand2_x0
xsubckt_1019_nand4_x0 2 1 1567 1571 1572 1593 1596 nand4_x0
xsubckt_339_nand3_x0 2 1 542 708 835 31 nand3_x0
xsubckt_1298_mx2_x2 1 1866 2 904 1344 50 mx2_x2
xsubckt_1764_sff1_x4 2 210 1 1953 114 sff1_x4
xsubckt_754_ao22_x2 1 1768 2 710 542 657 ao22_x2
xsubckt_680_nand3_x0 2 1 1838 263 269 141 nand3_x0
xsubckt_312_a4_x2 1 572 2 573 578 588 592 a4_x2
xsubckt_270_ao22_x2 1 614 2 736 732 628 ao22_x2
xsubckt_516_oa22_x2 1 367 2 368 390 797 oa22_x2
xsubckt_1374_nand2_x0 2 1 1275 580 150 nand2_x0
xsubckt_1523_ao22_x2 1 1132 2 803 1200 1243 ao22_x2
xsubckt_1799_sff1_x4 2 210 1 1925 37 sff1_x4
xsubckt_196_nand4_x0 2 1 695 23 834 26 836 nand4_x0
xsubckt_372_a4_x2 1 509 2 511 534 545 571 a4_x2
xsubckt_616_a4_x2 1 272 2 478 525 539 541 a4_x2
xsubckt_639_nand3_x0 2 1 249 543 719 43 nand3_x0
xsubckt_1284_nand2_x0 2 1 1356 1357 1362 nand2_x0
xsubckt_1455_o2_x2 1 1199 2 1200 802 o2_x2
xsubckt_1623_nand3_x0 2 1 1032 1181 1186 91 nand3_x0
xsubckt_980_nand3_x0 2 1 1602 1614 614 621 nand3_x0
xsubckt_908_oa22_x2 1 1636 2 1638 1640 890 oa22_x2
xsubckt_871_a4_x2 1 1668 2 784 788 795 909 a4_x2
xsubckt_853_nand2_x0 2 1 1682 1707 171 nand2_x0
xsubckt_820_oa22_x2 1 1971 2 1799 1792 1710 oa22_x2
xsubckt_283_nand2_x0 2 1 601 602 603 nand2_x0
xsubckt_420_a3_x2 2 462 1 621 729 766 a3_x2
xsubckt_1470_ao22_x2 1 1184 2 715 695 514 ao22_x2
xsubckt_1716_oa22_x2 1 939 2 1090 1075 1072 oa22_x2
xsubckt_1049_nand4_x0 2 1 1546 1581 612 650 753 nand4_x0
xsubckt_313_a2_x2 1 571 2 572 581 a2_x2
xsubckt_303_a2_x2 1 581 2 582 584 a2_x2
xsubckt_228_nand4_x0 2 1 659 662 708 26 836 nand4_x0
xsubckt_135_ao22_x2 1 769 2 71 89 774 ao22_x2
xsubckt_371_oa22_x2 1 510 2 12 653 513 oa22_x2
xsubckt_490_a3_x2 2 392 1 394 403 406 a3_x2
xsubckt_1406_nand2_x0 2 1 1246 1379 53 nand2_x0
xsubckt_1140_oa22_x2 1 1476 2 444 1478 1480 oa22_x2
xsubckt_816_oa22_x2 1 1713 2 1770 1771 849 oa22_x2
xsubckt_794_a3_x2 2 1732 1 1733 1736 1737 a3_x2
xsubckt_669_nand3_x0 2 1 222 263 269 142 nand3_x0
xsubckt_168_a2_x2 1 733 2 734 774 a2_x2
xsubckt_373_a2_x2 1 508 2 509 516 a2_x2
xsubckt_383_a2_x2 1 498 2 499 501 a2_x2
xsubckt_589_a3_x2 2 297 1 415 555 673 a3_x2
xsubckt_617_a2_x2 1 271 2 272 274 a2_x2
xsubckt_1427_ao22_x2 1 1227 2 1772 672 35 ao22_x2
xfeed_109 2 1 decap_w0
xfeed_108 2 1 decap_w0
xfeed_107 2 1 tie
xfeed_106 2 1 decap_w0
xfeed_105 2 1 decap_w0
xfeed_104 2 1 decap_w0
xfeed_103 2 1 tie
xfeed_102 2 1 decap_w0
xfeed_101 2 1 decap_w0
xfeed_100 2 1 decap_w0
xsubckt_973_nand2_x0 2 1 1607 647 38 nand2_x0
xsubckt_763_oa22_x2 1 1984 2 257 1792 1760 oa22_x2
xsubckt_724_oa22_x2 1 1797 2 249 550 881 oa22_x2
xsubckt_352_nand3_x0 2 1 529 658 680 794 nand3_x0
xsubckt_442_nand3_x0 2 1 440 449 640 693 nand3_x0
xsubckt_527_ao22_x2 1 356 2 448 441 357 ao22_x2
xsubckt_166_o2_x2 1 735 2 86 71 o2_x2
xsubckt_341_o2_x2 1 540 2 541 797 o2_x2
xsubckt_348_nand4_x0 2 1 533 658 680 831 27 nand4_x0
xsubckt_489_nand3_x0 2 1 393 645 769 771 nand3_x0
xsubckt_1364_a4_x2 1 1284 2 1285 1286 1287 550 a4_x2
xsubckt_1731_ao22_x2 1 924 2 925 926 949 ao22_x2
xsubckt_1880_sff1_x4 2 202 1 1853 156 sff1_x4
xfeed_119 2 1 decap_w0
xfeed_118 2 1 decap_w0
xfeed_117 2 1 decap_w0
xfeed_116 2 1 decap_w0
xfeed_115 2 1 tie
xfeed_114 2 1 tie
xfeed_113 2 1 tie
xfeed_112 2 1 tie
xfeed_111 2 1 tie
xfeed_110 2 1 tie
xsubckt_759_oa22_x2 1 1763 2 536 657 809 oa22_x2
xsubckt_236_oa22_x2 1 651 2 911 653 670 oa22_x2
xsubckt_511_nand4_x0 2 1 372 742 747 755 760 nand4_x0
xsubckt_525_nand2_x0 2 1 358 360 361 nand2_x0
xsubckt_1802_sff1_x4 2 205 1 1922 63 sff1_x4
xsubckt_1841_sff1_x4 2 209 1 1891 83 sff1_x4
xsubckt_1081_a2_x2 1 1520 2 1578 650 a2_x2
xsubckt_1071_a2_x2 1 1529 2 1530 1579 a2_x2
xsubckt_789_nand3_x0 2 1 1737 1767 1775 49 nand3_x0
xsubckt_675_o2_x2 1 216 2 256 862 o2_x2
xsubckt_255_mx2_x2 1 629 2 71 87 74 mx2_x2
xsubckt_1335_a2_x2 1 1310 2 1311 1312 a2_x2
xsubckt_1510_a2_x2 1 1145 2 1146 1227 a2_x2
xsubckt_1520_a2_x2 1 1135 2 1136 1154 a2_x2
xsubckt_1837_sff1_x4 2 211 1 1895 75 sff1_x4
xsubckt_1876_sff1_x4 2 207 1 1857 55 sff1_x4
xfeed_129 2 1 decap_w0
xfeed_128 2 1 decap_w0
xfeed_127 2 1 tie
xfeed_126 2 1 decap_w0
xfeed_125 2 1 decap_w0
xfeed_124 2 1 decap_w0
xfeed_123 2 1 decap_w0
xfeed_122 2 1 decap_w0
xfeed_121 2 1 tie
xfeed_120 2 1 tie
xsubckt_1149_mx2_x2 1 1890 2 1471 1469 102 mx2_x2
xsubckt_1148_mx2_x2 1 1469 2 586 1470 90 mx2_x2
xsubckt_1147_mx2_x2 1 1470 2 909 150 898 mx2_x2
xsubckt_1146_mx2_x2 1 1471 2 777 1472 585 mx2_x2
xsubckt_667_oa22_x2 1 189 2 288 229 224 oa22_x2
xsubckt_204_nand3_x0 2 1 687 784 23 834 nand3_x0
xsubckt_331_nand4_x0 2 1 553 691 795 833 20 nand4_x0
xsubckt_345_nand2_x0 2 1 536 543 713 nand2_x0
xsubckt_1355_a2_x2 1 1292 2 1293 1298 a2_x2
xsubckt_1365_a2_x2 1 1283 2 1284 1288 a2_x2
xsubckt_1436_oa22_x2 1 1218 2 1219 1221 40 oa22_x2
xsubckt_1629_a2_x2 1 1026 2 1027 1174 a2_x2
xsubckt_772_nand3_x0 2 1 1752 1767 1775 51 nand3_x0
xsubckt_292_nand3_x0 2 1 592 595 681 17 nand3_x0
xsubckt_378_nand4_x0 2 1 503 612 617 645 753 nand4_x0
xsubckt_1466_nand2_x0 2 1 1188 1190 1192 nand2_x0
xsubckt_1689_a2_x2 1 966 2 967 1212 a2_x2
xsubckt_1740_nxr2_x1 920 2 1 938 941 nxr2_x1
xsubckt_1784_sff1_x4 2 207 1 1939 124 sff1_x4
xfeed_139 2 1 decap_w0
xfeed_138 2 1 tie
xfeed_137 2 1 tie
xfeed_136 2 1 tie
xfeed_135 2 1 decap_w0
xfeed_134 2 1 decap_w0
xfeed_133 2 1 decap_w0
xfeed_132 2 1 decap_w0
xfeed_131 2 1 decap_w0
xfeed_130 2 1 decap_w0
xsubckt_1162_nor4_x0 2 1 1457 146 147 148 149 nor4_x0
xsubckt_682_nand3_x0 2 1 1836 263 268 125 nand3_x0
xsubckt_631_nand4_x0 2 1 257 258 259 260 261 nand4_x0
xsubckt_1305_oa22_x2 1 1337 2 49 1377 1339 oa22_x2
xsubckt_1490_o3_x2 1 1164 2 1167 1168 289 o3_x2
xsubckt_1582_ao22_x2 1 1073 2 1084 1086 1164 ao22_x2
xcmpt_abc_11873_new_n445_hfns_4 2 1 796 791 buf_x4
xcmpt_abc_11873_new_n445_hfns_3 2 1 791 792 buf_x4
xcmpt_abc_11873_new_n445_hfns_2 2 1 791 793 buf_x4
xcmpt_abc_11873_new_n445_hfns_1 2 1 791 794 buf_x4
xcmpt_abc_11873_new_n445_hfns_0 2 1 791 795 buf_x4
xcmpt_abc_11873_new_n443_hfns_2 2 1 801 798 buf_x4
xcmpt_abc_11873_new_n443_hfns_1 2 1 798 799 buf_x4
xcmpt_abc_11873_new_n443_hfns_0 2 1 798 800 buf_x4
xsubckt_1108_nand2_x0 2 1 1497 1498 1500 nand2_x0
xsubckt_678_nand4_x0 2 1 1839 1840 215 216 217 nand4_x0
xsubckt_1617_o2_x2 1 1038 2 1040 1042 o2_x2
xfeed_149 2 1 decap_w0
xfeed_148 2 1 decap_w0
xfeed_147 2 1 decap_w0
xfeed_146 2 1 tie
xfeed_145 2 1 tie
xfeed_144 2 1 decap_w0
xfeed_143 2 1 decap_w0
xfeed_142 2 1 decap_w0
xfeed_141 2 1 decap_w0
xfeed_140 2 1 decap_w0
xcmpt_abc_11873_new_n449_hfns_2 2 1 781 778 buf_x4
xcmpt_abc_11873_new_n449_hfns_1 2 1 778 779 buf_x4
xcmpt_abc_11873_new_n449_hfns_0 2 1 778 780 buf_x4
xcmpt_abc_11873_new_n448_hfns_2 2 1 785 782 buf_x4
xcmpt_abc_11873_new_n448_hfns_1 2 1 782 783 buf_x4
xcmpt_abc_11873_new_n448_hfns_0 2 1 782 784 buf_x4
xcmpt_abc_11873_new_n447_hfns_2 2 1 789 786 buf_x4
xcmpt_abc_11873_new_n447_hfns_1 2 1 786 787 buf_x4
xcmpt_abc_11873_new_n447_hfns_0 2 1 786 788 buf_x4
xsubckt_1145_nor3_x0 2 1 1472 38 109 42 nor3_x0
xsubckt_1018_nand2_x0 2 1 1568 648 869 nand2_x0
xsubckt_855_nand2_x0 2 1 1680 1780 88 nand2_x0
xsubckt_208_ao22_x2 1 683 2 687 710 12 ao22_x2
xsubckt_173_a3_x2 2 728 1 730 747 760 a3_x2
xsubckt_361_nand4_x0 2 1 520 658 679 17 832 nand4_x0
xsubckt_407_a3_x2 2 474 1 480 17 832 a3_x2
xsubckt_612_a3_x2 2 276 1 277 280 446 a3_x2
xsubckt_1578_ao22_x2 1 1077 2 1078 1087 1226 ao22_x2
xsubckt_261_a2_x2 1 623 2 624 774 a2_x2
xsubckt_487_a3_x2 2 395 1 396 397 398 a3_x2
xsubckt_505_a2_x2 1 378 2 742 747 a2_x2
xsubckt_624_nand3_x0 2 1 264 266 276 282 nand3_x0
xsubckt_1287_oa22_x2 1 1353 2 1373 1364 1356 oa22_x2
xsubckt_1408_nand2_x0 2 1 1244 580 147 nand2_x0
xsubckt_1486_ao22_x2 1 1168 2 1772 672 61 ao22_x2
xsubckt_1616_nor2_x0 2 1 1039 1040 1042 nor2_x0
xfeed_159 2 1 tie
xfeed_158 2 1 tie
xfeed_157 2 1 decap_w0
xfeed_156 2 1 decap_w0
xfeed_155 2 1 tie
xfeed_154 2 1 decap_w0
xfeed_153 2 1 decap_w0
xfeed_152 2 1 decap_w0
xfeed_151 2 1 decap_w0
xfeed_150 2 1 tie
xsubckt_1160_oa22_x2 1 1459 2 597 718 42 oa22_x2
xsubckt_1001_nand2_x0 2 1 1584 620 730 nand2_x0
xsubckt_692_a3_x2 2 1827 1 263 268 124 a3_x2
xsubckt_661_nand4_x0 2 1 229 231 232 233 234 nand4_x0
xsubckt_309_nxr2_x1 575 2 1 113 155 nxr2_x1
xsubckt_497_a3_x2 2 386 1 387 389 459 a3_x2
xsubckt_535_a2_x2 1 348 2 349 351 a2_x2
xsubckt_565_a2_x2 1 319 2 320 321 a2_x2
xsubckt_975_nand2_x0 2 1 1927 1606 1607 nand2_x0
xsubckt_783_oa22_x2 1 1742 2 536 657 806 oa22_x2
xsubckt_1591_oa22_x2 1 1064 2 150 1201 1066 oa22_x2
xfeed_209 2 1 tie
xfeed_208 2 1 decap_w0
xfeed_207 2 1 decap_w0
xfeed_206 2 1 decap_w0
xfeed_205 2 1 decap_w0
xfeed_204 2 1 decap_w0
xfeed_203 2 1 decap_w0
xfeed_202 2 1 tie
xfeed_201 2 1 decap_w0
xfeed_200 2 1 decap_w0
xfeed_169 2 1 decap_w0
xfeed_168 2 1 tie
xfeed_167 2 1 tie
xfeed_166 2 1 tie
xfeed_165 2 1 decap_w0
xfeed_164 2 1 decap_w0
xfeed_163 2 1 decap_w0
xfeed_162 2 1 decap_w0
xfeed_161 2 1 tie
xfeed_160 2 1 decap_w0
xsubckt_834_nand3_x0 2 1 1698 1767 1775 57 nand3_x0
xsubckt_104_mx2_x2 1 809 2 903 823 824 mx2_x2
xsubckt_1301_nand2_x0 2 1 1341 1343 550 nand2_x0
xsubckt_1552_oa22_x2 1 1103 2 148 1201 1105 oa22_x2
xsubckt_795_nand2_x0 2 1 1974 1732 1738 nand2_x0
xsubckt_779_oa22_x2 1 1976 2 229 1792 1746 oa22_x2
xsubckt_691_oa22_x2 1 187 2 288 1833 1828 oa22_x2
xsubckt_652_oa22_x2 1 237 2 253 700 896 oa22_x2
xsubckt_106_mx2_x2 1 808 2 904 820 821 mx2_x2
xsubckt_108_mx2_x2 1 807 2 904 817 818 mx2_x2
xsubckt_1822_sff1_x4 2 211 1 93 101 sff1_x4
xsubckt_1861_sff1_x4 2 206 1 1872 171 sff1_x4
xfeed_219 2 1 tie
xfeed_218 2 1 decap_w0
xfeed_217 2 1 decap_w0
xfeed_216 2 1 decap_w0
xfeed_215 2 1 tie
xfeed_214 2 1 decap_w0
xfeed_213 2 1 decap_w0
xfeed_212 2 1 decap_w0
xfeed_211 2 1 decap_w0
xfeed_210 2 1 decap_w0
xfeed_179 2 1 decap_w0
xfeed_178 2 1 decap_w0
xfeed_177 2 1 decap_w0
xfeed_176 2 1 decap_w0
xfeed_175 2 1 decap_w0
xfeed_174 2 1 tie
xfeed_173 2 1 decap_w0
xfeed_172 2 1 tie
xfeed_171 2 1 decap_w0
xfeed_170 2 1 tie
xsubckt_1213_a2_x2 1 1409 2 594 657 a2_x2
xsubckt_1099_oa22_x2 1 1903 2 41 777 4 oa22_x2
xsubckt_398_o2_x2 1 483 2 484 797 o2_x2
xsubckt_564_nand3_x0 2 1 320 597 719 800 nand3_x0
xsubckt_1385_nand3_x0 2 1 1265 591 792 172 nand3_x0
xsubckt_1479_a3_x2 2 1175 1 1177 1190 1192 a3_x2
xsubckt_1509_oa22_x2 1 1146 2 257 1205 1147 oa22_x2
xsubckt_1818_sff1_x4 2 209 1 1906 33 sff1_x4
xsubckt_1857_sff1_x4 2 206 1 1876 175 sff1_x4
xsubckt_1078_nand2_x0 2 1 1523 647 826 nand2_x0
xsubckt_827_nand2_x0 2 1 1970 1704 1709 nand2_x0
xsubckt_474_nand3_x0 2 1 408 610 740 767 nand3_x0
xsubckt_600_nand2_x0 2 1 287 707 715 nand2_x0
xsubckt_1348_mx2_x2 1 1861 2 904 1299 45 mx2_x2
xsubckt_1694_ao22_x2 1 961 2 964 965 969 ao22_x2
xsubckt_1722_a2_x2 1 933 2 1120 1136 a2_x2
xsubckt_1736_mx2_x2 1 1851 2 904 921 153 mx2_x2
xsubckt_1737_mx2_x2 1 1850 2 904 947 152 mx2_x2
xsubckt_1738_mx2_x2 1 1849 2 904 945 151 mx2_x2
xsubckt_1739_mx2_x2 1 1848 2 904 951 150 mx2_x2
xfeed_229 2 1 decap_w0
xfeed_228 2 1 tie
xfeed_227 2 1 tie
xfeed_226 2 1 decap_w0
xfeed_225 2 1 decap_w0
xfeed_224 2 1 decap_w0
xfeed_223 2 1 tie
xfeed_222 2 1 tie
xfeed_221 2 1 decap_w0
xfeed_220 2 1 decap_w0
xfeed_189 2 1 decap_w0
xfeed_188 2 1 decap_w0
xfeed_187 2 1 tie
xfeed_186 2 1 decap_w0
xfeed_185 2 1 decap_w0
xfeed_184 2 1 decap_w0
xfeed_183 2 1 tie
xfeed_182 2 1 decap_w0
xfeed_181 2 1 tie
xfeed_180 2 1 decap_w0
xsubckt_864_nand3_x0 2 1 1673 1767 1775 52 nand3_x0
xsubckt_257_nand2_x0 2 1 627 629 774 nand2_x0
xsubckt_167_nand2_x0 2 1 734 843 71 nand2_x0
xsubckt_510_nand2_x0 2 1 373 437 454 nand2_x0
xsubckt_1558_nand2_x0 2 1 1097 1098 1099 nand2_x0
xsubckt_1577_a2_x2 1 1078 2 1079 1174 a2_x2
xsubckt_1595_nand3_x0 2 1 1060 1181 1186 90 nand3_x0
xsubckt_1655_ao22_x2 1 1000 2 1004 1006 1189 ao22_x2
xsubckt_1765_sff1_x4 2 205 1 183 32 sff1_x4
xsubckt_1325_oa22_x2 1 1319 2 47 1377 1321 oa22_x2
xsubckt_1698_mx2_x2 1 957 2 992 989 990 mx2_x2
xfeed_239 2 1 decap_w0
xfeed_238 2 1 tie
xfeed_237 2 1 decap_w0
xfeed_236 2 1 decap_w0
xfeed_235 2 1 decap_w0
xfeed_234 2 1 decap_w0
xfeed_233 2 1 decap_w0
xfeed_232 2 1 tie
xfeed_231 2 1 decap_w0
xfeed_230 2 1 decap_w0
xfeed_199 2 1 decap_w0
xfeed_198 2 1 decap_w0
xfeed_197 2 1 decap_w0
xfeed_196 2 1 decap_w0
xfeed_195 2 1 decap_w0
xfeed_194 2 1 decap_w0
xfeed_193 2 1 decap_w0
xfeed_192 2 1 tie
xfeed_191 2 1 decap_w0
xfeed_190 2 1 decap_w0
xsubckt_909_nxr2_x1 1635 2 1 1637 148 nxr2_x1
xsubckt_240_nand2_x0 2 1 644 650 900 nand2_x0
xsubckt_237_a4_x2 1 650 2 784 788 795 9 a4_x2
xsubckt_227_a4_x2 1 660 2 662 708 26 836 a4_x2
xsubckt_1094_nand4_x0 2 1 1509 1600 621 742 747 nand4_x0
xsubckt_984_nand3_x0 2 1 1599 627 731 734 nand3_x0
xsubckt_857_nand2_x0 2 1 1979 1679 1683 nand2_x0
xsubckt_806_nand3_x0 2 1 1722 1767 1775 47 nand3_x0
xsubckt_150_nand2_x0 2 1 754 757 759 nand2_x0
xsubckt_326_nand3_x0 2 1 558 570 681 717 nand3_x0
xfeed_249 2 1 decap_w0
xfeed_248 2 1 decap_w0
xfeed_247 2 1 tie
xfeed_246 2 1 decap_w0
xfeed_245 2 1 tie
xfeed_244 2 1 decap_w0
xfeed_243 2 1 decap_w0
xfeed_242 2 1 decap_w0
xfeed_241 2 1 decap_w0
xfeed_240 2 1 decap_w0
xfeed_0 2 1 decap_w0
xsubckt_1220_nand3_x0 2 1 1402 1418 1783 287 nand3_x0
xsubckt_991_a4_x2 1 1594 2 628 729 742 747 a4_x2
xsubckt_197_nand2_x0 2 1 694 698 713 nand2_x0
xsubckt_365_a3_x2 2 516 1 517 523 531 a3_x2
xsubckt_540_a3_x2 2 343 1 344 523 531 a3_x2
xsubckt_1664_nxr2_x1 991 2 1 1002 1164 nxr2_x1
xfeed_9 2 1 decap_w0
xfeed_8 2 1 decap_w0
xfeed_7 2 1 tie
xfeed_6 2 1 decap_w0
xfeed_5 2 1 decap_w0
xfeed_4 2 1 tie
xfeed_3 2 1 decap_w0
xfeed_2 2 1 decap_w0
xfeed_1 2 1 decap_w0
xsubckt_1180_oa22_x2 1 1442 2 493 687 710 oa22_x2
xsubckt_1141_oa22_x2 1 1475 2 1477 1479 917 oa22_x2
xsubckt_1130_nand3_x0 2 1 1485 1486 1668 899 nand3_x0
xsubckt_844_a3_x2 2 1689 1 1690 1691 1692 a3_x2
xsubckt_453_a2_x2 1 429 2 430 432 a2_x2
xfeed_259 2 1 decap_w0
xfeed_258 2 1 decap_w0
xfeed_257 2 1 tie
xfeed_256 2 1 tie
xfeed_255 2 1 decap_w0
xfeed_254 2 1 tie
xfeed_253 2 1 tie
xfeed_252 2 1 decap_w0
xfeed_251 2 1 decap_w0
xfeed_250 2 1 decap_w0
xsubckt_1091_nand2_x0 2 1 1511 1512 1617 nand2_x0
xsubckt_305_nand4_x0 2 1 579 691 794 23 834 nand4_x0
xsubckt_298_a2_x2 1 586 2 597 718 a2_x2
xsubckt_285_o4_x2 1 599 2 601 636 641 651 o4_x2
xsubckt_280_oa22_x2 1 604 2 645 607 632 oa22_x2
xsubckt_446_nand3_x0 2 1 436 438 741 747 nand3_x0
xsubckt_746_nand3_x0 2 1 1776 1777 1779 1781 nand3_x0
xsubckt_725_oa22_x2 1 1796 2 253 700 887 oa22_x2
xsubckt_209_nor2_x0 2 1 682 4 9 nor2_x0
xsubckt_528_ao22_x2 1 355 2 736 732 627 ao22_x2
xsubckt_1340_nand3_x0 2 1 1306 591 793 176 nand3_x0
xsubckt_1414_a4_x2 1 1238 2 1239 1251 1260 1269 a4_x2
xsubckt_1533_oa22_x2 1 1122 2 1125 1126 1175 oa22_x2
xfeed_309 2 1 decap_w0
xfeed_308 2 1 decap_w0
xfeed_307 2 1 decap_w0
xfeed_306 2 1 decap_w0
xfeed_305 2 1 decap_w0
xfeed_304 2 1 decap_w0
xfeed_303 2 1 decap_w0
xfeed_302 2 1 decap_w0
xfeed_301 2 1 decap_w0
xfeed_300 2 1 decap_w0
xfeed_269 2 1 decap_w0
xfeed_268 2 1 decap_w0
xfeed_267 2 1 decap_w0
xfeed_266 2 1 decap_w0
xfeed_265 2 1 tie
xfeed_264 2 1 tie
xfeed_263 2 1 decap_w0
xfeed_262 2 1 decap_w0
xfeed_261 2 1 decap_w0
xfeed_260 2 1 decap_w0
xsubckt_1123_nand2_x0 2 1 1492 672 112 nand2_x0
xsubckt_1111_a2_x2 1 1495 2 398 518 a2_x2
xsubckt_799_oa22_x2 1 1728 2 536 657 804 oa22_x2
xsubckt_656_nand3_x0 2 1 234 262 268 119 nand3_x0
xsubckt_1512_a3_x2 2 1143 1 698 793 47 a3_x2
xsubckt_1803_sff1_x4 2 205 1 1921 62 sff1_x4
xsubckt_1842_sff1_x4 2 210 1 1890 102 sff1_x4
xsubckt_1881_sff1_x4 2 202 1 1852 155 sff1_x4
xsubckt_1205_ao22_x2 1 1417 2 497 698 792 ao22_x2
xsubckt_515_nand4_x0 2 1 368 369 374 383 386 nand4_x0
xsubckt_1283_ao22_x2 1 1357 2 893 1385 1358 ao22_x2
xsubckt_1367_a3_x2 2 1281 1 1282 1291 1300 a3_x2
xsubckt_1529_oa22_x2 1 1126 2 1140 1142 1188 oa22_x2
xsubckt_1600_a2_x2 1 1055 2 1056 1174 a2_x2
xsubckt_1610_a2_x2 1 1045 2 1049 1053 a2_x2
xsubckt_1877_sff1_x4 2 207 1 1856 54 sff1_x4
xfeed_319 2 1 decap_w0
xfeed_318 2 1 decap_w0
xfeed_317 2 1 decap_w0
xfeed_316 2 1 decap_w0
xfeed_315 2 1 decap_w0
xfeed_314 2 1 decap_w0
xfeed_313 2 1 decap_w0
xfeed_312 2 1 decap_w0
xfeed_311 2 1 decap_w0
xfeed_310 2 1 decap_w0
xfeed_279 2 1 decap_w0
xfeed_278 2 1 tie
xfeed_277 2 1 decap_w0
xfeed_276 2 1 tie
xfeed_275 2 1 tie
xfeed_274 2 1 decap_w0
xfeed_273 2 1 decap_w0
xfeed_272 2 1 tie
xfeed_271 2 1 tie
xfeed_270 2 1 decap_w0
xsubckt_1156_mx2_x2 1 1462 2 1463 86 146 mx2_x2
xsubckt_1070_nand3_x0 2 1 1530 1600 620 761 nand3_x0
xsubckt_1011_o3_x2 1 1574 2 1576 1582 1588 o3_x2
xsubckt_829_nand2_x0 2 1 1702 1707 175 nand2_x0
xsubckt_349_nand2_x0 2 1 532 754 761 nand2_x0
xsubckt_386_nand3_x0 2 1 495 497 680 718 nand3_x0
xsubckt_602_nand2_x0 2 1 285 286 14 nand2_x0
xsubckt_1465_a2_x2 1 1189 2 1190 1192 a2_x2
xsubckt_1476_oa22_x2 1 1178 2 1180 1187 1188 oa22_x2
xsubckt_1719_a2_x2 1 936 2 1093 1110 a2_x2
xsubckt_1750_sff1_x4 2 208 1 1967 144 sff1_x4
xsubckt_1838_sff1_x4 2 211 1 1894 74 sff1_x4
xsubckt_1157_mx2_x2 1 1889 2 1464 66 1462 mx2_x2
xsubckt_1152_ao22_x2 1 1466 2 263 268 67 ao22_x2
xsubckt_740_ao22_x2 1 1782 2 719 713 497 ao22_x2
xsubckt_296_nand3_x0 2 1 588 591 713 800 nand3_x0
xsubckt_169_nand2_x0 2 1 732 734 774 nand2_x0
xsubckt_1437_oa22_x2 1 1217 2 577 686 889 oa22_x2
xsubckt_1785_sff1_x4 2 206 1 1938 123 sff1_x4
xfeed_329 2 1 decap_w0
xfeed_328 2 1 decap_w0
xfeed_327 2 1 decap_w0
xfeed_326 2 1 decap_w0
xfeed_325 2 1 decap_w0
xfeed_324 2 1 decap_w0
xfeed_323 2 1 decap_w0
xfeed_322 2 1 decap_w0
xfeed_321 2 1 decap_w0
xfeed_320 2 1 decap_w0
xfeed_289 2 1 decap_w0
xfeed_288 2 1 decap_w0
xfeed_287 2 1 decap_w0
xfeed_286 2 1 decap_w0
xfeed_285 2 1 decap_w0
xfeed_284 2 1 decap_w0
xfeed_283 2 1 decap_w0
xfeed_282 2 1 decap_w0
xfeed_281 2 1 decap_w0
xfeed_280 2 1 decap_w0
xsubckt_1228_o2_x2 1 1394 2 1395 1399 o2_x2
xsubckt_1153_nand2_x0 2 1 1465 1668 906 nand2_x0
xsubckt_1163_nor4_x0 2 1 1456 150 151 152 153 nor4_x0
xsubckt_990_nand2_x0 2 1 1595 648 870 nand2_x0
xsubckt_812_nand2_x0 2 1 1972 1717 1723 nand2_x0
xsubckt_203_a3_x2 2 688 1 784 23 834 a3_x2
xsubckt_330_a4_x2 1 554 2 691 795 833 20 a4_x2
xsubckt_332_nand2_x0 2 1 552 554 681 nand2_x0
xsubckt_455_nand4_x0 2 1 427 610 645 740 766 nand4_x0
xsubckt_1505_ao22_x2 1 1150 2 1203 1789 153 ao22_x2
xsubckt_1670_nand3_x0 2 1 985 698 795 59 nand3_x0
xfeed_339 2 1 decap_w0
xfeed_338 2 1 decap_w0
xfeed_337 2 1 decap_w0
xfeed_336 2 1 decap_w0
xfeed_335 2 1 decap_w0
xfeed_334 2 1 decap_w0
xfeed_333 2 1 decap_w0
xfeed_332 2 1 decap_w0
xfeed_331 2 1 decap_w0
xfeed_330 2 1 decap_w0
xfeed_299 2 1 decap_w0
xfeed_298 2 1 decap_w0
xfeed_297 2 1 decap_w0
xfeed_296 2 1 decap_w0
xfeed_295 2 1 decap_w0
xfeed_294 2 1 decap_w0
xfeed_293 2 1 decap_w0
xfeed_292 2 1 decap_w0
xfeed_291 2 1 decap_w0
xfeed_290 2 1 decap_w0
xspare_buffer_19 2 1 7 3 buf_x4
xspare_buffer_18 2 1 212 200 buf_x4
xspare_buffer_17 2 1 212 201 buf_x4
xspare_buffer_16 2 1 212 202 buf_x4
xspare_buffer_15 2 1 7 4 buf_x4
xspare_buffer_14 2 1 212 203 buf_x4
xspare_buffer_13 2 1 212 204 buf_x4
xspare_buffer_12 2 1 212 205 buf_x4
xspare_buffer_11 2 1 7 5 buf_x4
xspare_buffer_10 2 1 212 206 buf_x4
xsubckt_859_nand2_x0 2 1 1677 1707 170 nand2_x0
xsubckt_195_a4_x2 1 699 2 23 834 26 836 a4_x2
xsubckt_152_nand2_x0 2 1 752 755 760 nand2_x0
xsubckt_328_nand3_x0 2 1 556 566 717 800 nand3_x0
xsubckt_379_nand2_x0 2 1 502 698 795 nand2_x0
xsubckt_1402_nand3_x0 2 1 1249 1251 1260 1269 nand3_x0
xsubckt_1453_nand2_x0 2 1 1201 1204 1790 nand2_x0
xsubckt_1017_ao22_x2 1 1922 2 1570 1573 1595 ao22_x2
xsubckt_732_a3_x2 2 1790 1 1791 559 583 a3_x2
xsubckt_718_nand3_x0 2 1 1803 262 269 130 nand3_x0
xsubckt_684_a4_x2 1 1834 2 1835 1836 1837 1838 a4_x2
xsubckt_321_a2_x2 1 563 2 566 713 a2_x2
xsubckt_557_a3_x2 2 327 1 328 335 338 a3_x2
xsubckt_628_nand3_x0 2 1 260 262 268 121 nand3_x0
xsubckt_1363_nand2_x0 2 1 1285 580 151 nand2_x0
xfeed_349 2 1 decap_w0
xfeed_348 2 1 decap_w0
xfeed_347 2 1 decap_w0
xfeed_346 2 1 decap_w0
xfeed_345 2 1 decap_w0
xfeed_344 2 1 decap_w0
xfeed_343 2 1 decap_w0
xfeed_342 2 1 decap_w0
xfeed_341 2 1 decap_w0
xfeed_340 2 1 decap_w0
xsubckt_1183_nand2_x0 2 1 1439 1442 1443 nand2_x0
xsubckt_810_a2_x2 1 1718 2 1719 1720 a2_x2
xsubckt_752_a3_x2 2 1770 1 579 656 694 a3_x2
xsubckt_311_nand3_x0 2 1 573 574 591 794 nand3_x0
xsubckt_362_nand2_x0 2 1 519 528 16 nand2_x0
xsubckt_538_nand3_x0 2 1 345 679 688 713 nand3_x0
xsubckt_615_a2_x2 1 273 2 478 541 a2_x2
xsubckt_1179_nand3_x0 2 1 1443 783 793 23 nand3_x0
xsubckt_979_nand2_x0 2 1 1603 647 37 nand2_x0
xsubckt_870_a2_x2 1 1841 2 159 102 a2_x2
xsubckt_842_nand2_x0 2 1 1691 1780 90 nand2_x0
xsubckt_448_nand3_x0 2 1 434 437 613 645 nand3_x0
xsubckt_499_nand2_x0 2 1 384 385 608 nand2_x0
xsubckt_1573_nand2_x0 2 1 1082 1083 1085 nand2_x0
xfeed_359 2 1 tie
xfeed_358 2 1 decap_w0
xfeed_357 2 1 decap_w0
xfeed_356 2 1 decap_w0
xfeed_355 2 1 decap_w0
xfeed_354 2 1 decap_w0
xfeed_353 2 1 decap_w0
xfeed_352 2 1 decap_w0
xfeed_351 2 1 decap_w0
xfeed_350 2 1 decap_w0
xsubckt_959_a2_x2 1 1617 2 504 650 a2_x2
xsubckt_268_nand3_x0 2 1 616 620 729 766 nand3_x0
xsubckt_182_nand2_x0 2 1 715 831 27 nand2_x0
xsubckt_110_mx2_x2 1 806 2 903 814 815 mx2_x2
xsubckt_509_ao22_x2 1 374 2 436 381 375 ao22_x2
xsubckt_1342_a4_x2 1 1304 2 1305 1306 1307 550 a4_x2
xsubckt_1252_nand3_x0 2 1 1386 1783 593 709 nand3_x0
xsubckt_658_nand3_x0 2 1 232 262 269 135 nand3_x0
xsubckt_178_nand3_x0 2 1 723 788 26 836 nand3_x0
xsubckt_112_mx2_x2 1 805 2 903 811 812 mx2_x2
xsubckt_114_mx2_x2 1 804 2 904 838 839 mx2_x2
xsubckt_116_mx2_x2 1 803 2 904 841 842 mx2_x2
xsubckt_633_o2_x2 1 255 2 256 865 o2_x2
xsubckt_1393_nand2_x0 2 1 1258 1379 54 nand2_x0
xsubckt_1713_ao22_x2 1 942 2 952 1045 1046 ao22_x2
xsubckt_1823_sff1_x4 2 211 1 92 100 sff1_x4
xsubckt_1862_sff1_x4 2 206 1 1871 170 sff1_x4
.ends arlet6502_cts_r
