* Coriolis Structural SPICE Driver
* Generated on Apr 11, 2023, 23:42
* Cell/Subckt "Arlet6502".
* 
* INTERF vss
* INTERF vdd
* INTERF reset
* INTERF clk
* INTERF WE
* INTERF RDY
* INTERF NMI
* INTERF IRQ
* INTERF DO[7]
* INTERF DO[6]
* INTERF DO[5]
* INTERF DO[4]
* INTERF DO[3]
* INTERF DO[2]
* INTERF DO[1]
* INTERF DO[0]
* INTERF DI[7]
* INTERF DI[6]
* INTERF DI[5]
* INTERF DI[4]
* INTERF DI[3]
* INTERF DI[2]
* INTERF DI[1]
* INTERF DI[0]
* INTERF A[9]
* INTERF A[8]
* INTERF A[7]
* INTERF A[6]
* INTERF A[5]
* INTERF A[4]
* INTERF A[3]
* INTERF A[2]
* INTERF A[15]
* INTERF A[14]
* INTERF A[13]
* INTERF A[12]
* INTERF A[11]
* INTERF A[10]
* INTERF A[1]
* INTERF A[0]

* Terminal models (aka standard cells) used througout all the hierarchy.
.include mx2_x2.spi
.include a3_x2.spi
.include oa22_x2.spi
.include ao22_x2.spi
.include o2_x2.spi
.include nand3_x0.spi
.include nand2_x0.spi
.include sff1_x4.spi
.include a2_x2.spi
.include nand4_x0.spi
.include o4_x2.spi
.include nxr2_x1.spi
.include a4_x2.spi
.include nor2_x0.spi
.include mx3_x2.spi
.include inv_x0.spi
.include nor3_x0.spi
.include nor4_x0.spi
.include o3_x2.spi
.include xr2_x1.spi

* Non-terminal models (part of the user's design hierarchy).

.subckt Arlet6502 0 1 2 9 1720 1721 1722 1874 1875 1876 1877 1878 1879 1880 1881 1882 1883 1884 1885 1886 1887 1888 1889 1890 1891 1892 1893 1894 1895 1896 1897 1898 1899 1900 1901 1902 1903 1904 1905 1906
* NET     0 = vss
* NET     1 = vdd
* NET     2 = reset
* NET     3 = flatten_MOS6502_auto_fsm_map_cc_288_map_fsm_1405_Y[5]
* NET     4 = flatten_MOS6502_auto_fsm_map_cc_288_map_fsm_1405_Y[4]
* NET     5 = flatten_MOS6502_auto_fsm_map_cc_288_map_fsm_1405_Y[3]
* NET     6 = flatten_MOS6502_auto_fsm_map_cc_288_map_fsm_1405_Y[2]
* NET     7 = flatten_MOS6502_auto_fsm_map_cc_288_map_fsm_1405_Y[1]
* NET     8 = flatten_MOS6502_auto_fsm_map_cc_288_map_fsm_1405_Y[0]
* NET     9 = clk
* NET    10 = abc_11873_new_n999
* NET    11 = abc_11873_new_n998
* NET    12 = abc_11873_new_n997
* NET    13 = abc_11873_new_n996
* NET    14 = abc_11873_new_n995
* NET    15 = abc_11873_new_n994
* NET    16 = abc_11873_new_n993
* NET    17 = abc_11873_new_n992
* NET    18 = abc_11873_new_n991
* NET    19 = abc_11873_new_n989
* NET    20 = abc_11873_new_n988
* NET    21 = abc_11873_new_n987
* NET    22 = abc_11873_new_n986
* NET    23 = abc_11873_new_n985
* NET    24 = abc_11873_new_n984
* NET    25 = abc_11873_new_n983
* NET    26 = abc_11873_new_n982
* NET    27 = abc_11873_new_n981
* NET    28 = abc_11873_new_n980
* NET    29 = abc_11873_new_n979
* NET    30 = abc_11873_new_n977
* NET    31 = abc_11873_new_n976
* NET    32 = abc_11873_new_n975
* NET    33 = abc_11873_new_n974
* NET    34 = abc_11873_new_n973
* NET    35 = abc_11873_new_n972
* NET    36 = abc_11873_new_n971
* NET    37 = abc_11873_new_n970
* NET    38 = abc_11873_new_n969
* NET    39 = abc_11873_new_n968
* NET    40 = abc_11873_new_n967
* NET    41 = abc_11873_new_n965
* NET    42 = abc_11873_new_n964
* NET    43 = abc_11873_new_n963
* NET    44 = abc_11873_new_n962
* NET    45 = abc_11873_new_n961
* NET    46 = abc_11873_new_n960
* NET    47 = abc_11873_new_n959
* NET    48 = abc_11873_new_n958
* NET    49 = abc_11873_new_n957
* NET    50 = abc_11873_new_n956
* NET    51 = abc_11873_new_n955
* NET    52 = abc_11873_new_n954
* NET    53 = abc_11873_new_n953
* NET    54 = abc_11873_new_n952
* NET    55 = abc_11873_new_n951
* NET    56 = abc_11873_new_n950
* NET    57 = abc_11873_new_n949
* NET    58 = abc_11873_new_n948
* NET    59 = abc_11873_new_n947
* NET    60 = abc_11873_new_n946
* NET    61 = abc_11873_new_n945
* NET    62 = abc_11873_new_n944
* NET    63 = abc_11873_new_n943
* NET    64 = abc_11873_new_n942
* NET    65 = abc_11873_new_n941
* NET    66 = abc_11873_new_n940
* NET    67 = abc_11873_new_n939
* NET    68 = abc_11873_new_n938
* NET    69 = abc_11873_new_n937
* NET    70 = abc_11873_new_n936
* NET    71 = abc_11873_new_n935
* NET    72 = abc_11873_new_n934
* NET    73 = abc_11873_new_n933
* NET    74 = abc_11873_new_n932
* NET    75 = abc_11873_new_n931
* NET    76 = abc_11873_new_n930
* NET    77 = abc_11873_new_n929
* NET    78 = abc_11873_new_n928
* NET    79 = abc_11873_new_n927
* NET    80 = abc_11873_new_n925
* NET    81 = abc_11873_new_n924
* NET    82 = abc_11873_new_n923
* NET    83 = abc_11873_new_n922
* NET    84 = abc_11873_new_n921
* NET    85 = abc_11873_new_n920
* NET    86 = abc_11873_new_n918
* NET    87 = abc_11873_new_n917
* NET    88 = abc_11873_new_n916
* NET    89 = abc_11873_new_n915
* NET    90 = abc_11873_new_n914
* NET    91 = abc_11873_new_n913
* NET    92 = abc_11873_new_n912
* NET    93 = abc_11873_new_n911
* NET    94 = abc_11873_new_n910
* NET    95 = abc_11873_new_n909
* NET    96 = abc_11873_new_n908
* NET    97 = abc_11873_new_n906
* NET    98 = abc_11873_new_n905
* NET    99 = abc_11873_new_n904
* NET   100 = abc_11873_new_n903
* NET   101 = abc_11873_new_n902
* NET   102 = abc_11873_new_n901
* NET   103 = abc_11873_new_n900
* NET   104 = abc_11873_new_n899
* NET   105 = abc_11873_new_n897
* NET   106 = abc_11873_new_n896
* NET   107 = abc_11873_new_n895
* NET   108 = abc_11873_new_n894
* NET   109 = abc_11873_new_n893
* NET   110 = abc_11873_new_n892
* NET   111 = abc_11873_new_n891
* NET   112 = abc_11873_new_n890
* NET   113 = abc_11873_new_n889
* NET   114 = abc_11873_new_n888
* NET   115 = abc_11873_new_n887
* NET   116 = abc_11873_new_n886
* NET   117 = abc_11873_new_n885
* NET   118 = abc_11873_new_n884
* NET   119 = abc_11873_new_n883
* NET   120 = abc_11873_new_n882
* NET   121 = abc_11873_new_n881
* NET   122 = abc_11873_new_n880
* NET   123 = abc_11873_new_n879
* NET   124 = abc_11873_new_n878
* NET   125 = abc_11873_new_n877
* NET   126 = abc_11873_new_n876
* NET   127 = abc_11873_new_n875
* NET   128 = abc_11873_new_n874
* NET   129 = abc_11873_new_n873
* NET   130 = abc_11873_new_n872
* NET   131 = abc_11873_new_n871
* NET   132 = abc_11873_new_n870
* NET   133 = abc_11873_new_n869
* NET   134 = abc_11873_new_n868
* NET   135 = abc_11873_new_n866
* NET   136 = abc_11873_new_n865
* NET   137 = abc_11873_new_n864
* NET   138 = abc_11873_new_n863
* NET   139 = abc_11873_new_n862
* NET   140 = abc_11873_new_n861
* NET   141 = abc_11873_new_n860
* NET   142 = abc_11873_new_n859
* NET   143 = abc_11873_new_n858
* NET   144 = abc_11873_new_n857
* NET   145 = abc_11873_new_n856
* NET   146 = abc_11873_new_n855
* NET   147 = abc_11873_new_n854
* NET   148 = abc_11873_new_n853
* NET   149 = abc_11873_new_n852
* NET   150 = abc_11873_new_n851
* NET   151 = abc_11873_new_n850
* NET   152 = abc_11873_new_n849
* NET   153 = abc_11873_new_n848
* NET   154 = abc_11873_new_n847
* NET   155 = abc_11873_new_n846
* NET   156 = abc_11873_new_n845
* NET   157 = abc_11873_new_n844
* NET   158 = abc_11873_new_n843
* NET   159 = abc_11873_new_n842
* NET   160 = abc_11873_new_n841
* NET   161 = abc_11873_new_n840
* NET   162 = abc_11873_new_n839
* NET   163 = abc_11873_new_n838
* NET   164 = abc_11873_new_n837
* NET   165 = abc_11873_new_n836
* NET   166 = abc_11873_new_n835
* NET   167 = abc_11873_new_n834
* NET   168 = abc_11873_new_n833
* NET   169 = abc_11873_new_n832
* NET   170 = abc_11873_new_n831
* NET   171 = abc_11873_new_n830
* NET   172 = abc_11873_new_n829
* NET   173 = abc_11873_new_n828
* NET   174 = abc_11873_new_n827
* NET   175 = abc_11873_new_n826
* NET   176 = abc_11873_new_n825
* NET   177 = abc_11873_new_n824
* NET   178 = abc_11873_new_n823
* NET   179 = abc_11873_new_n822
* NET   180 = abc_11873_new_n821
* NET   181 = abc_11873_new_n820
* NET   182 = abc_11873_new_n819
* NET   183 = abc_11873_new_n818
* NET   184 = abc_11873_new_n817
* NET   185 = abc_11873_new_n816
* NET   186 = abc_11873_new_n814
* NET   187 = abc_11873_new_n813
* NET   188 = abc_11873_new_n812
* NET   189 = abc_11873_new_n811
* NET   190 = abc_11873_new_n810
* NET   191 = abc_11873_new_n809
* NET   192 = abc_11873_new_n808
* NET   193 = abc_11873_new_n807
* NET   194 = abc_11873_new_n806
* NET   195 = abc_11873_new_n805
* NET   196 = abc_11873_new_n804
* NET   197 = abc_11873_new_n803
* NET   198 = abc_11873_new_n802
* NET   199 = abc_11873_new_n801
* NET   200 = abc_11873_new_n800
* NET   201 = abc_11873_new_n799
* NET   202 = abc_11873_new_n798
* NET   203 = abc_11873_new_n797
* NET   204 = abc_11873_new_n796
* NET   205 = abc_11873_new_n795
* NET   206 = abc_11873_new_n794
* NET   207 = abc_11873_new_n793
* NET   208 = abc_11873_new_n792
* NET   209 = abc_11873_new_n791
* NET   210 = abc_11873_new_n790
* NET   211 = abc_11873_new_n789
* NET   212 = abc_11873_new_n788
* NET   213 = abc_11873_new_n787
* NET   214 = abc_11873_new_n786
* NET   215 = abc_11873_new_n785
* NET   216 = abc_11873_new_n784
* NET   217 = abc_11873_new_n783
* NET   218 = abc_11873_new_n782
* NET   219 = abc_11873_new_n781
* NET   220 = abc_11873_new_n780
* NET   221 = abc_11873_new_n779
* NET   222 = abc_11873_new_n778
* NET   223 = abc_11873_new_n777
* NET   224 = abc_11873_new_n776
* NET   225 = abc_11873_new_n775
* NET   226 = abc_11873_new_n774
* NET   227 = abc_11873_new_n773
* NET   228 = abc_11873_new_n772
* NET   229 = abc_11873_new_n771
* NET   230 = abc_11873_new_n770
* NET   231 = abc_11873_new_n769
* NET   232 = abc_11873_new_n768
* NET   233 = abc_11873_new_n767
* NET   234 = abc_11873_new_n766
* NET   235 = abc_11873_new_n765
* NET   236 = abc_11873_new_n764
* NET   237 = abc_11873_new_n763
* NET   238 = abc_11873_new_n762
* NET   239 = abc_11873_new_n761
* NET   240 = abc_11873_new_n760
* NET   241 = abc_11873_new_n759
* NET   242 = abc_11873_new_n758
* NET   243 = abc_11873_new_n757
* NET   244 = abc_11873_new_n756
* NET   245 = abc_11873_new_n755
* NET   246 = abc_11873_new_n754
* NET   247 = abc_11873_new_n753
* NET   248 = abc_11873_new_n752
* NET   249 = abc_11873_new_n751
* NET   250 = abc_11873_new_n750
* NET   251 = abc_11873_new_n749
* NET   252 = abc_11873_new_n748
* NET   253 = abc_11873_new_n747
* NET   254 = abc_11873_new_n746
* NET   255 = abc_11873_new_n745
* NET   256 = abc_11873_new_n744
* NET   257 = abc_11873_new_n743
* NET   258 = abc_11873_new_n742
* NET   259 = abc_11873_new_n740
* NET   260 = abc_11873_new_n739
* NET   261 = abc_11873_new_n738
* NET   262 = abc_11873_new_n737
* NET   263 = abc_11873_new_n736
* NET   264 = abc_11873_new_n735
* NET   265 = abc_11873_new_n734
* NET   266 = abc_11873_new_n733
* NET   267 = abc_11873_new_n732
* NET   268 = abc_11873_new_n731
* NET   269 = abc_11873_new_n730
* NET   270 = abc_11873_new_n729
* NET   271 = abc_11873_new_n728
* NET   272 = abc_11873_new_n727
* NET   273 = abc_11873_new_n726
* NET   274 = abc_11873_new_n725
* NET   275 = abc_11873_new_n724
* NET   276 = abc_11873_new_n723
* NET   277 = abc_11873_new_n722
* NET   278 = abc_11873_new_n721
* NET   279 = abc_11873_new_n720
* NET   280 = abc_11873_new_n719
* NET   281 = abc_11873_new_n718
* NET   282 = abc_11873_new_n717
* NET   283 = abc_11873_new_n716
* NET   284 = abc_11873_new_n715
* NET   285 = abc_11873_new_n714
* NET   286 = abc_11873_new_n713
* NET   287 = abc_11873_new_n712
* NET   288 = abc_11873_new_n711
* NET   289 = abc_11873_new_n710
* NET   290 = abc_11873_new_n709
* NET   291 = abc_11873_new_n708
* NET   292 = abc_11873_new_n707
* NET   293 = abc_11873_new_n706
* NET   294 = abc_11873_new_n705
* NET   295 = abc_11873_new_n704
* NET   296 = abc_11873_new_n703
* NET   297 = abc_11873_new_n702
* NET   298 = abc_11873_new_n701
* NET   299 = abc_11873_new_n700
* NET   300 = abc_11873_new_n699
* NET   301 = abc_11873_new_n698
* NET   302 = abc_11873_new_n697
* NET   303 = abc_11873_new_n696
* NET   304 = abc_11873_new_n695
* NET   305 = abc_11873_new_n694
* NET   306 = abc_11873_new_n693
* NET   307 = abc_11873_new_n692
* NET   308 = abc_11873_new_n691
* NET   309 = abc_11873_new_n690
* NET   310 = abc_11873_new_n689
* NET   311 = abc_11873_new_n688
* NET   312 = abc_11873_new_n687
* NET   313 = abc_11873_new_n686
* NET   314 = abc_11873_new_n685
* NET   315 = abc_11873_new_n684
* NET   316 = abc_11873_new_n683
* NET   317 = abc_11873_new_n682
* NET   318 = abc_11873_new_n681
* NET   319 = abc_11873_new_n680
* NET   320 = abc_11873_new_n679
* NET   321 = abc_11873_new_n678
* NET   322 = abc_11873_new_n677
* NET   323 = abc_11873_new_n676
* NET   324 = abc_11873_new_n675
* NET   325 = abc_11873_new_n674
* NET   326 = abc_11873_new_n673
* NET   327 = abc_11873_new_n672
* NET   328 = abc_11873_new_n671
* NET   329 = abc_11873_new_n670
* NET   330 = abc_11873_new_n669
* NET   331 = abc_11873_new_n668
* NET   332 = abc_11873_new_n667
* NET   333 = abc_11873_new_n666
* NET   334 = abc_11873_new_n665
* NET   335 = abc_11873_new_n664
* NET   336 = abc_11873_new_n663
* NET   337 = abc_11873_new_n662
* NET   338 = abc_11873_new_n661
* NET   339 = abc_11873_new_n660
* NET   340 = abc_11873_new_n659
* NET   341 = abc_11873_new_n658
* NET   342 = abc_11873_new_n657
* NET   343 = abc_11873_new_n656
* NET   344 = abc_11873_new_n655
* NET   345 = abc_11873_new_n654
* NET   346 = abc_11873_new_n653
* NET   347 = abc_11873_new_n652
* NET   348 = abc_11873_new_n651
* NET   349 = abc_11873_new_n650
* NET   350 = abc_11873_new_n649
* NET   351 = abc_11873_new_n648
* NET   352 = abc_11873_new_n647
* NET   353 = abc_11873_new_n646
* NET   354 = abc_11873_new_n645
* NET   355 = abc_11873_new_n644
* NET   356 = abc_11873_new_n643
* NET   357 = abc_11873_new_n642
* NET   358 = abc_11873_new_n641
* NET   359 = abc_11873_new_n640
* NET   360 = abc_11873_new_n639
* NET   361 = abc_11873_new_n638
* NET   362 = abc_11873_new_n637
* NET   363 = abc_11873_new_n636
* NET   364 = abc_11873_new_n635
* NET   365 = abc_11873_new_n634
* NET   366 = abc_11873_new_n633
* NET   367 = abc_11873_new_n632
* NET   368 = abc_11873_new_n631
* NET   369 = abc_11873_new_n630
* NET   370 = abc_11873_new_n629
* NET   371 = abc_11873_new_n628
* NET   372 = abc_11873_new_n627
* NET   373 = abc_11873_new_n626
* NET   374 = abc_11873_new_n625
* NET   375 = abc_11873_new_n624
* NET   376 = abc_11873_new_n623
* NET   377 = abc_11873_new_n622
* NET   378 = abc_11873_new_n621
* NET   379 = abc_11873_new_n620
* NET   380 = abc_11873_new_n619
* NET   381 = abc_11873_new_n618
* NET   382 = abc_11873_new_n617
* NET   383 = abc_11873_new_n616
* NET   384 = abc_11873_new_n615
* NET   385 = abc_11873_new_n614
* NET   386 = abc_11873_new_n613
* NET   387 = abc_11873_new_n612
* NET   388 = abc_11873_new_n611
* NET   389 = abc_11873_new_n610
* NET   390 = abc_11873_new_n609
* NET   391 = abc_11873_new_n608
* NET   392 = abc_11873_new_n607
* NET   393 = abc_11873_new_n606
* NET   394 = abc_11873_new_n605
* NET   395 = abc_11873_new_n604
* NET   396 = abc_11873_new_n603
* NET   397 = abc_11873_new_n602
* NET   398 = abc_11873_new_n601
* NET   399 = abc_11873_new_n600
* NET   400 = abc_11873_new_n599
* NET   401 = abc_11873_new_n598
* NET   402 = abc_11873_new_n597
* NET   403 = abc_11873_new_n596
* NET   404 = abc_11873_new_n595
* NET   405 = abc_11873_new_n594
* NET   406 = abc_11873_new_n593
* NET   407 = abc_11873_new_n592
* NET   408 = abc_11873_new_n591
* NET   409 = abc_11873_new_n590
* NET   410 = abc_11873_new_n589
* NET   411 = abc_11873_new_n588
* NET   412 = abc_11873_new_n587
* NET   413 = abc_11873_new_n586
* NET   414 = abc_11873_new_n585
* NET   415 = abc_11873_new_n584
* NET   416 = abc_11873_new_n583
* NET   417 = abc_11873_new_n582
* NET   418 = abc_11873_new_n581
* NET   419 = abc_11873_new_n580
* NET   420 = abc_11873_new_n579
* NET   421 = abc_11873_new_n578
* NET   422 = abc_11873_new_n577
* NET   423 = abc_11873_new_n576
* NET   424 = abc_11873_new_n575
* NET   425 = abc_11873_new_n574
* NET   426 = abc_11873_new_n573
* NET   427 = abc_11873_new_n572
* NET   428 = abc_11873_new_n571
* NET   429 = abc_11873_new_n570
* NET   430 = abc_11873_new_n569
* NET   431 = abc_11873_new_n568
* NET   432 = abc_11873_new_n567
* NET   433 = abc_11873_new_n566
* NET   434 = abc_11873_new_n565
* NET   435 = abc_11873_new_n564
* NET   436 = abc_11873_new_n563
* NET   437 = abc_11873_new_n562
* NET   438 = abc_11873_new_n561
* NET   439 = abc_11873_new_n560
* NET   440 = abc_11873_new_n559
* NET   441 = abc_11873_new_n558
* NET   442 = abc_11873_new_n557
* NET   443 = abc_11873_new_n556
* NET   444 = abc_11873_new_n555
* NET   445 = abc_11873_new_n554
* NET   446 = abc_11873_new_n553
* NET   447 = abc_11873_new_n552
* NET   448 = abc_11873_new_n551
* NET   449 = abc_11873_new_n550
* NET   450 = abc_11873_new_n549
* NET   451 = abc_11873_new_n548
* NET   452 = abc_11873_new_n547
* NET   453 = abc_11873_new_n546
* NET   454 = abc_11873_new_n545
* NET   455 = abc_11873_new_n544
* NET   456 = abc_11873_new_n543
* NET   457 = abc_11873_new_n542
* NET   458 = abc_11873_new_n541
* NET   459 = abc_11873_new_n540
* NET   460 = abc_11873_new_n539
* NET   461 = abc_11873_new_n538
* NET   462 = abc_11873_new_n537
* NET   463 = abc_11873_new_n536
* NET   464 = abc_11873_new_n535
* NET   465 = abc_11873_new_n534
* NET   466 = abc_11873_new_n533
* NET   467 = abc_11873_new_n532
* NET   468 = abc_11873_new_n531
* NET   469 = abc_11873_new_n530
* NET   470 = abc_11873_new_n529
* NET   471 = abc_11873_new_n528
* NET   472 = abc_11873_new_n527
* NET   473 = abc_11873_new_n526
* NET   474 = abc_11873_new_n525
* NET   475 = abc_11873_new_n524
* NET   476 = abc_11873_new_n523
* NET   477 = abc_11873_new_n522
* NET   478 = abc_11873_new_n521
* NET   479 = abc_11873_new_n520
* NET   480 = abc_11873_new_n519
* NET   481 = abc_11873_new_n518
* NET   482 = abc_11873_new_n517
* NET   483 = abc_11873_new_n516
* NET   484 = abc_11873_new_n515
* NET   485 = abc_11873_new_n514
* NET   486 = abc_11873_new_n513
* NET   487 = abc_11873_new_n512
* NET   488 = abc_11873_new_n511
* NET   489 = abc_11873_new_n510
* NET   490 = abc_11873_new_n509
* NET   491 = abc_11873_new_n508
* NET   492 = abc_11873_new_n507
* NET   493 = abc_11873_new_n506
* NET   494 = abc_11873_new_n505
* NET   495 = abc_11873_new_n504
* NET   496 = abc_11873_new_n503
* NET   497 = abc_11873_new_n502
* NET   498 = abc_11873_new_n501
* NET   499 = abc_11873_new_n500
* NET   500 = abc_11873_new_n499
* NET   501 = abc_11873_new_n498
* NET   502 = abc_11873_new_n497
* NET   503 = abc_11873_new_n496
* NET   504 = abc_11873_new_n495
* NET   505 = abc_11873_new_n494
* NET   506 = abc_11873_new_n493
* NET   507 = abc_11873_new_n492
* NET   508 = abc_11873_new_n491
* NET   509 = abc_11873_new_n490
* NET   510 = abc_11873_new_n489
* NET   511 = abc_11873_new_n488
* NET   512 = abc_11873_new_n487
* NET   513 = abc_11873_new_n486
* NET   514 = abc_11873_new_n485
* NET   515 = abc_11873_new_n484
* NET   516 = abc_11873_new_n483
* NET   517 = abc_11873_new_n482
* NET   518 = abc_11873_new_n481
* NET   519 = abc_11873_new_n480
* NET   520 = abc_11873_new_n479
* NET   521 = abc_11873_new_n478
* NET   522 = abc_11873_new_n477
* NET   523 = abc_11873_new_n476
* NET   524 = abc_11873_new_n475
* NET   525 = abc_11873_new_n474
* NET   526 = abc_11873_new_n473
* NET   527 = abc_11873_new_n472
* NET   528 = abc_11873_new_n471
* NET   529 = abc_11873_new_n470
* NET   530 = abc_11873_new_n469
* NET   531 = abc_11873_new_n468
* NET   532 = abc_11873_new_n467
* NET   533 = abc_11873_new_n466
* NET   534 = abc_11873_new_n465
* NET   535 = abc_11873_new_n464
* NET   536 = abc_11873_new_n463
* NET   537 = abc_11873_new_n462
* NET   538 = abc_11873_new_n461
* NET   539 = abc_11873_new_n460
* NET   540 = abc_11873_new_n459
* NET   541 = abc_11873_new_n458
* NET   542 = abc_11873_new_n457
* NET   543 = abc_11873_new_n456
* NET   544 = abc_11873_new_n455
* NET   545 = abc_11873_new_n454
* NET   546 = abc_11873_new_n453
* NET   547 = abc_11873_new_n452
* NET   548 = abc_11873_new_n451
* NET   549 = abc_11873_new_n450
* NET   550 = abc_11873_new_n449
* NET   551 = abc_11873_new_n448
* NET   552 = abc_11873_new_n447
* NET   553 = abc_11873_new_n446
* NET   554 = abc_11873_new_n445
* NET   555 = abc_11873_new_n444
* NET   556 = abc_11873_new_n443
* NET   557 = abc_11873_new_n441
* NET   558 = abc_11873_new_n439
* NET   559 = abc_11873_new_n437
* NET   560 = abc_11873_new_n435
* NET   561 = abc_11873_new_n433
* NET   562 = abc_11873_new_n431
* NET   563 = abc_11873_new_n429
* NET   564 = abc_11873_new_n427
* NET   565 = abc_11873_new_n426
* NET   566 = abc_11873_new_n425
* NET   567 = abc_11873_new_n424
* NET   568 = abc_11873_new_n423
* NET   569 = abc_11873_new_n422
* NET   570 = abc_11873_new_n421
* NET   571 = abc_11873_new_n420
* NET   572 = abc_11873_new_n419
* NET   573 = abc_11873_new_n418
* NET   574 = abc_11873_new_n417
* NET   575 = abc_11873_new_n416
* NET   576 = abc_11873_new_n415
* NET   577 = abc_11873_new_n414
* NET   578 = abc_11873_new_n413
* NET   579 = abc_11873_new_n412
* NET   580 = abc_11873_new_n411
* NET   581 = abc_11873_new_n410
* NET   582 = abc_11873_new_n409
* NET   583 = abc_11873_new_n408
* NET   584 = abc_11873_new_n407
* NET   585 = abc_11873_new_n406
* NET   586 = abc_11873_new_n405
* NET   587 = abc_11873_new_n404
* NET   588 = abc_11873_new_n403
* NET   589 = abc_11873_new_n402
* NET   590 = abc_11873_new_n401
* NET   591 = abc_11873_new_n400
* NET   592 = abc_11873_new_n399
* NET   593 = abc_11873_new_n398
* NET   594 = abc_11873_new_n397
* NET   595 = abc_11873_new_n396
* NET   596 = abc_11873_new_n395
* NET   597 = abc_11873_new_n394
* NET   598 = abc_11873_new_n393
* NET   599 = abc_11873_new_n392
* NET   600 = abc_11873_new_n391
* NET   601 = abc_11873_new_n390
* NET   602 = abc_11873_new_n389
* NET   603 = abc_11873_new_n388
* NET   604 = abc_11873_new_n387
* NET   605 = abc_11873_new_n386
* NET   606 = abc_11873_new_n385
* NET   607 = abc_11873_new_n384
* NET   608 = abc_11873_new_n383
* NET   609 = abc_11873_new_n382
* NET   610 = abc_11873_new_n381
* NET   611 = abc_11873_new_n380
* NET   612 = abc_11873_new_n379
* NET   613 = abc_11873_new_n378
* NET   614 = abc_11873_new_n377
* NET   615 = abc_11873_new_n376
* NET   616 = abc_11873_new_n375
* NET   617 = abc_11873_new_n374
* NET   618 = abc_11873_new_n373
* NET   619 = abc_11873_new_n372
* NET   620 = abc_11873_new_n371
* NET   621 = abc_11873_new_n370
* NET   622 = abc_11873_new_n369
* NET   623 = abc_11873_new_n368
* NET   624 = abc_11873_new_n367
* NET   625 = abc_11873_new_n366
* NET   626 = abc_11873_new_n365
* NET   627 = abc_11873_new_n364
* NET   628 = abc_11873_new_n363
* NET   629 = abc_11873_new_n362
* NET   630 = abc_11873_new_n361
* NET   631 = abc_11873_new_n360
* NET   632 = abc_11873_new_n359
* NET   633 = abc_11873_new_n358
* NET   634 = abc_11873_new_n357
* NET   635 = abc_11873_new_n356
* NET   636 = abc_11873_new_n355
* NET   637 = abc_11873_new_n354
* NET   638 = abc_11873_new_n353
* NET   639 = abc_11873_new_n352
* NET   640 = abc_11873_new_n351
* NET   641 = abc_11873_new_n350
* NET   642 = abc_11873_new_n349
* NET   643 = abc_11873_new_n348
* NET   644 = abc_11873_new_n347
* NET   645 = abc_11873_new_n346
* NET   646 = abc_11873_new_n345
* NET   647 = abc_11873_new_n344
* NET   648 = abc_11873_new_n343
* NET   649 = abc_11873_new_n342
* NET   650 = abc_11873_new_n341
* NET   651 = abc_11873_new_n340
* NET   652 = abc_11873_new_n339
* NET   653 = abc_11873_new_n338
* NET   654 = abc_11873_new_n337
* NET   655 = abc_11873_new_n336
* NET   656 = abc_11873_new_n335
* NET   657 = abc_11873_new_n334
* NET   658 = abc_11873_new_n333
* NET   659 = abc_11873_new_n332
* NET   660 = abc_11873_new_n331
* NET   661 = abc_11873_new_n330
* NET   662 = abc_11873_new_n329
* NET   663 = abc_11873_new_n328
* NET   664 = abc_11873_new_n327
* NET   665 = abc_11873_new_n326
* NET   666 = abc_11873_new_n325
* NET   667 = abc_11873_new_n324
* NET   668 = abc_11873_new_n323
* NET   669 = abc_11873_new_n2069
* NET   670 = abc_11873_new_n2068
* NET   671 = abc_11873_new_n2063
* NET   672 = abc_11873_new_n2058
* NET   673 = abc_11873_new_n2057
* NET   674 = abc_11873_new_n2055
* NET   675 = abc_11873_new_n2054
* NET   676 = abc_11873_new_n2053
* NET   677 = abc_11873_new_n2052
* NET   678 = abc_11873_new_n2051
* NET   679 = abc_11873_new_n2050
* NET   680 = abc_11873_new_n2049
* NET   681 = abc_11873_new_n2048
* NET   682 = abc_11873_new_n2047
* NET   683 = abc_11873_new_n2046
* NET   684 = abc_11873_new_n2045
* NET   685 = abc_11873_new_n2044
* NET   686 = abc_11873_new_n2043
* NET   687 = abc_11873_new_n2042
* NET   688 = abc_11873_new_n2041
* NET   689 = abc_11873_new_n2040
* NET   690 = abc_11873_new_n2039
* NET   691 = abc_11873_new_n2038
* NET   692 = abc_11873_new_n2037
* NET   693 = abc_11873_new_n2036
* NET   694 = abc_11873_new_n2035
* NET   695 = abc_11873_new_n2034
* NET   696 = abc_11873_new_n2033
* NET   697 = abc_11873_new_n2032
* NET   698 = abc_11873_new_n2031
* NET   699 = abc_11873_new_n2030
* NET   700 = abc_11873_new_n2029
* NET   701 = abc_11873_new_n2028
* NET   702 = abc_11873_new_n2027
* NET   703 = abc_11873_new_n2026
* NET   704 = abc_11873_new_n2025
* NET   705 = abc_11873_new_n2024
* NET   706 = abc_11873_new_n2023
* NET   707 = abc_11873_new_n2022
* NET   708 = abc_11873_new_n2021
* NET   709 = abc_11873_new_n2020
* NET   710 = abc_11873_new_n2019
* NET   711 = abc_11873_new_n2018
* NET   712 = abc_11873_new_n2017
* NET   713 = abc_11873_new_n2016
* NET   714 = abc_11873_new_n2015
* NET   715 = abc_11873_new_n2014
* NET   716 = abc_11873_new_n2013
* NET   717 = abc_11873_new_n2012
* NET   718 = abc_11873_new_n2011
* NET   719 = abc_11873_new_n2010
* NET   720 = abc_11873_new_n2009
* NET   721 = abc_11873_new_n2008
* NET   722 = abc_11873_new_n2007
* NET   723 = abc_11873_new_n2006
* NET   724 = abc_11873_new_n2005
* NET   725 = abc_11873_new_n2004
* NET   726 = abc_11873_new_n2003
* NET   727 = abc_11873_new_n2002
* NET   728 = abc_11873_new_n2001
* NET   729 = abc_11873_new_n2000
* NET   730 = abc_11873_new_n1999
* NET   731 = abc_11873_new_n1998
* NET   732 = abc_11873_new_n1997
* NET   733 = abc_11873_new_n1996
* NET   734 = abc_11873_new_n1995
* NET   735 = abc_11873_new_n1994
* NET   736 = abc_11873_new_n1993
* NET   737 = abc_11873_new_n1992
* NET   738 = abc_11873_new_n1991
* NET   739 = abc_11873_new_n1990
* NET   740 = abc_11873_new_n1989
* NET   741 = abc_11873_new_n1988
* NET   742 = abc_11873_new_n1987
* NET   743 = abc_11873_new_n1986
* NET   744 = abc_11873_new_n1985
* NET   745 = abc_11873_new_n1984
* NET   746 = abc_11873_new_n1983
* NET   747 = abc_11873_new_n1982
* NET   748 = abc_11873_new_n1981
* NET   749 = abc_11873_new_n1980
* NET   750 = abc_11873_new_n1979
* NET   751 = abc_11873_new_n1978
* NET   752 = abc_11873_new_n1977
* NET   753 = abc_11873_new_n1976
* NET   754 = abc_11873_new_n1975
* NET   755 = abc_11873_new_n1974
* NET   756 = abc_11873_new_n1973
* NET   757 = abc_11873_new_n1972
* NET   758 = abc_11873_new_n1971
* NET   759 = abc_11873_new_n1970
* NET   760 = abc_11873_new_n1969
* NET   761 = abc_11873_new_n1968
* NET   762 = abc_11873_new_n1967
* NET   763 = abc_11873_new_n1966
* NET   764 = abc_11873_new_n1965
* NET   765 = abc_11873_new_n1964
* NET   766 = abc_11873_new_n1963
* NET   767 = abc_11873_new_n1962
* NET   768 = abc_11873_new_n1961
* NET   769 = abc_11873_new_n1960
* NET   770 = abc_11873_new_n1959
* NET   771 = abc_11873_new_n1958
* NET   772 = abc_11873_new_n1957
* NET   773 = abc_11873_new_n1956
* NET   774 = abc_11873_new_n1955
* NET   775 = abc_11873_new_n1954
* NET   776 = abc_11873_new_n1953
* NET   777 = abc_11873_new_n1952
* NET   778 = abc_11873_new_n1951
* NET   779 = abc_11873_new_n1950
* NET   780 = abc_11873_new_n1949
* NET   781 = abc_11873_new_n1948
* NET   782 = abc_11873_new_n1947
* NET   783 = abc_11873_new_n1946
* NET   784 = abc_11873_new_n1945
* NET   785 = abc_11873_new_n1944
* NET   786 = abc_11873_new_n1943
* NET   787 = abc_11873_new_n1942
* NET   788 = abc_11873_new_n1941
* NET   789 = abc_11873_new_n1940
* NET   790 = abc_11873_new_n1939
* NET   791 = abc_11873_new_n1938
* NET   792 = abc_11873_new_n1937
* NET   793 = abc_11873_new_n1936
* NET   794 = abc_11873_new_n1935
* NET   795 = abc_11873_new_n1934
* NET   796 = abc_11873_new_n1933
* NET   797 = abc_11873_new_n1932
* NET   798 = abc_11873_new_n1931
* NET   799 = abc_11873_new_n1930
* NET   800 = abc_11873_new_n1929
* NET   801 = abc_11873_new_n1928
* NET   802 = abc_11873_new_n1927
* NET   803 = abc_11873_new_n1926
* NET   804 = abc_11873_new_n1925
* NET   805 = abc_11873_new_n1924
* NET   806 = abc_11873_new_n1923
* NET   807 = abc_11873_new_n1922
* NET   808 = abc_11873_new_n1921
* NET   809 = abc_11873_new_n1920
* NET   810 = abc_11873_new_n1919
* NET   811 = abc_11873_new_n1918
* NET   812 = abc_11873_new_n1917
* NET   813 = abc_11873_new_n1916
* NET   814 = abc_11873_new_n1915
* NET   815 = abc_11873_new_n1914
* NET   816 = abc_11873_new_n1913
* NET   817 = abc_11873_new_n1912
* NET   818 = abc_11873_new_n1911
* NET   819 = abc_11873_new_n1910
* NET   820 = abc_11873_new_n1909
* NET   821 = abc_11873_new_n1908
* NET   822 = abc_11873_new_n1907
* NET   823 = abc_11873_new_n1906
* NET   824 = abc_11873_new_n1905
* NET   825 = abc_11873_new_n1904
* NET   826 = abc_11873_new_n1903
* NET   827 = abc_11873_new_n1902
* NET   828 = abc_11873_new_n1901
* NET   829 = abc_11873_new_n1900
* NET   830 = abc_11873_new_n1899
* NET   831 = abc_11873_new_n1898
* NET   832 = abc_11873_new_n1897
* NET   833 = abc_11873_new_n1896
* NET   834 = abc_11873_new_n1895
* NET   835 = abc_11873_new_n1894
* NET   836 = abc_11873_new_n1893
* NET   837 = abc_11873_new_n1892
* NET   838 = abc_11873_new_n1891
* NET   839 = abc_11873_new_n1890
* NET   840 = abc_11873_new_n1889
* NET   841 = abc_11873_new_n1888
* NET   842 = abc_11873_new_n1887
* NET   843 = abc_11873_new_n1886
* NET   844 = abc_11873_new_n1885
* NET   845 = abc_11873_new_n1884
* NET   846 = abc_11873_new_n1883
* NET   847 = abc_11873_new_n1882
* NET   848 = abc_11873_new_n1881
* NET   849 = abc_11873_new_n1880
* NET   850 = abc_11873_new_n1879
* NET   851 = abc_11873_new_n1878
* NET   852 = abc_11873_new_n1877
* NET   853 = abc_11873_new_n1876
* NET   854 = abc_11873_new_n1875
* NET   855 = abc_11873_new_n1874
* NET   856 = abc_11873_new_n1873
* NET   857 = abc_11873_new_n1872
* NET   858 = abc_11873_new_n1871
* NET   859 = abc_11873_new_n1870
* NET   860 = abc_11873_new_n1869
* NET   861 = abc_11873_new_n1868
* NET   862 = abc_11873_new_n1867
* NET   863 = abc_11873_new_n1866
* NET   864 = abc_11873_new_n1865
* NET   865 = abc_11873_new_n1864
* NET   866 = abc_11873_new_n1863
* NET   867 = abc_11873_new_n1862
* NET   868 = abc_11873_new_n1861
* NET   869 = abc_11873_new_n1860
* NET   870 = abc_11873_new_n1859
* NET   871 = abc_11873_new_n1858
* NET   872 = abc_11873_new_n1857
* NET   873 = abc_11873_new_n1856
* NET   874 = abc_11873_new_n1855
* NET   875 = abc_11873_new_n1854
* NET   876 = abc_11873_new_n1853
* NET   877 = abc_11873_new_n1852
* NET   878 = abc_11873_new_n1851
* NET   879 = abc_11873_new_n1850
* NET   880 = abc_11873_new_n1849
* NET   881 = abc_11873_new_n1848
* NET   882 = abc_11873_new_n1847
* NET   883 = abc_11873_new_n1846
* NET   884 = abc_11873_new_n1845
* NET   885 = abc_11873_new_n1844
* NET   886 = abc_11873_new_n1843
* NET   887 = abc_11873_new_n1842
* NET   888 = abc_11873_new_n1841
* NET   889 = abc_11873_new_n1840
* NET   890 = abc_11873_new_n1839
* NET   891 = abc_11873_new_n1838
* NET   892 = abc_11873_new_n1837
* NET   893 = abc_11873_new_n1836
* NET   894 = abc_11873_new_n1835
* NET   895 = abc_11873_new_n1834
* NET   896 = abc_11873_new_n1833
* NET   897 = abc_11873_new_n1832
* NET   898 = abc_11873_new_n1831
* NET   899 = abc_11873_new_n1830
* NET   900 = abc_11873_new_n1829
* NET   901 = abc_11873_new_n1828
* NET   902 = abc_11873_new_n1827
* NET   903 = abc_11873_new_n1825
* NET   904 = abc_11873_new_n1824
* NET   905 = abc_11873_new_n1823
* NET   906 = abc_11873_new_n1822
* NET   907 = abc_11873_new_n1821
* NET   908 = abc_11873_new_n1820
* NET   909 = abc_11873_new_n1819
* NET   910 = abc_11873_new_n1818
* NET   911 = abc_11873_new_n1817
* NET   912 = abc_11873_new_n1816
* NET   913 = abc_11873_new_n1815
* NET   914 = abc_11873_new_n1814
* NET   915 = abc_11873_new_n1813
* NET   916 = abc_11873_new_n1812
* NET   917 = abc_11873_new_n1811
* NET   918 = abc_11873_new_n1810
* NET   919 = abc_11873_new_n1809
* NET   920 = abc_11873_new_n1808
* NET   921 = abc_11873_new_n1807
* NET   922 = abc_11873_new_n1806
* NET   923 = abc_11873_new_n1805
* NET   924 = abc_11873_new_n1804
* NET   925 = abc_11873_new_n1803
* NET   926 = abc_11873_new_n1802
* NET   927 = abc_11873_new_n1801
* NET   928 = abc_11873_new_n1800
* NET   929 = abc_11873_new_n1799
* NET   930 = abc_11873_new_n1798
* NET   931 = abc_11873_new_n1797
* NET   932 = abc_11873_new_n1796
* NET   933 = abc_11873_new_n1795
* NET   934 = abc_11873_new_n1794
* NET   935 = abc_11873_new_n1793
* NET   936 = abc_11873_new_n1792
* NET   937 = abc_11873_new_n1791
* NET   938 = abc_11873_new_n1790
* NET   939 = abc_11873_new_n1789
* NET   940 = abc_11873_new_n1788
* NET   941 = abc_11873_new_n1787
* NET   942 = abc_11873_new_n1786
* NET   943 = abc_11873_new_n1785
* NET   944 = abc_11873_new_n1784
* NET   945 = abc_11873_new_n1783
* NET   946 = abc_11873_new_n1782
* NET   947 = abc_11873_new_n1781
* NET   948 = abc_11873_new_n1780
* NET   949 = abc_11873_new_n1779
* NET   950 = abc_11873_new_n1778
* NET   951 = abc_11873_new_n1777
* NET   952 = abc_11873_new_n1776
* NET   953 = abc_11873_new_n1775
* NET   954 = abc_11873_new_n1774
* NET   955 = abc_11873_new_n1773
* NET   956 = abc_11873_new_n1772
* NET   957 = abc_11873_new_n1771
* NET   958 = abc_11873_new_n1770
* NET   959 = abc_11873_new_n1769
* NET   960 = abc_11873_new_n1768
* NET   961 = abc_11873_new_n1767
* NET   962 = abc_11873_new_n1766
* NET   963 = abc_11873_new_n1765
* NET   964 = abc_11873_new_n1764
* NET   965 = abc_11873_new_n1763
* NET   966 = abc_11873_new_n1762
* NET   967 = abc_11873_new_n1761
* NET   968 = abc_11873_new_n1760
* NET   969 = abc_11873_new_n1759
* NET   970 = abc_11873_new_n1758
* NET   971 = abc_11873_new_n1757
* NET   972 = abc_11873_new_n1756
* NET   973 = abc_11873_new_n1755
* NET   974 = abc_11873_new_n1754
* NET   975 = abc_11873_new_n1753
* NET   976 = abc_11873_new_n1752
* NET   977 = abc_11873_new_n1751
* NET   978 = abc_11873_new_n1750
* NET   979 = abc_11873_new_n1749
* NET   980 = abc_11873_new_n1747
* NET   981 = abc_11873_new_n1746
* NET   982 = abc_11873_new_n1745
* NET   983 = abc_11873_new_n1744
* NET   984 = abc_11873_new_n1743
* NET   985 = abc_11873_new_n1742
* NET   986 = abc_11873_new_n1741
* NET   987 = abc_11873_new_n1740
* NET   988 = abc_11873_new_n1738
* NET   989 = abc_11873_new_n1737
* NET   990 = abc_11873_new_n1736
* NET   991 = abc_11873_new_n1735
* NET   992 = abc_11873_new_n1734
* NET   993 = abc_11873_new_n1733
* NET   994 = abc_11873_new_n1732
* NET   995 = abc_11873_new_n1731
* NET   996 = abc_11873_new_n1730
* NET   997 = abc_11873_new_n1729
* NET   998 = abc_11873_new_n1727
* NET   999 = abc_11873_new_n1726
* NET  1000 = abc_11873_new_n1725
* NET  1001 = abc_11873_new_n1724
* NET  1002 = abc_11873_new_n1723
* NET  1003 = abc_11873_new_n1722
* NET  1004 = abc_11873_new_n1721
* NET  1005 = abc_11873_new_n1720
* NET  1006 = abc_11873_new_n1719
* NET  1007 = abc_11873_new_n1718
* NET  1008 = abc_11873_new_n1717
* NET  1009 = abc_11873_new_n1716
* NET  1010 = abc_11873_new_n1714
* NET  1011 = abc_11873_new_n1713
* NET  1012 = abc_11873_new_n1712
* NET  1013 = abc_11873_new_n1711
* NET  1014 = abc_11873_new_n1710
* NET  1015 = abc_11873_new_n1709
* NET  1016 = abc_11873_new_n1708
* NET  1017 = abc_11873_new_n1707
* NET  1018 = abc_11873_new_n1706
* NET  1019 = abc_11873_new_n1704
* NET  1020 = abc_11873_new_n1703
* NET  1021 = abc_11873_new_n1702
* NET  1022 = abc_11873_new_n1701
* NET  1023 = abc_11873_new_n1700
* NET  1024 = abc_11873_new_n1699
* NET  1025 = abc_11873_new_n1698
* NET  1026 = abc_11873_new_n1697
* NET  1027 = abc_11873_new_n1696
* NET  1028 = abc_11873_new_n1695
* NET  1029 = abc_11873_new_n1693
* NET  1030 = abc_11873_new_n1692
* NET  1031 = abc_11873_new_n1691
* NET  1032 = abc_11873_new_n1690
* NET  1033 = abc_11873_new_n1689
* NET  1034 = abc_11873_new_n1688
* NET  1035 = abc_11873_new_n1687
* NET  1036 = abc_11873_new_n1686
* NET  1037 = abc_11873_new_n1685
* NET  1038 = abc_11873_new_n1684
* NET  1039 = abc_11873_new_n1683
* NET  1040 = abc_11873_new_n1682
* NET  1041 = abc_11873_new_n1680
* NET  1042 = abc_11873_new_n1679
* NET  1043 = abc_11873_new_n1678
* NET  1044 = abc_11873_new_n1677
* NET  1045 = abc_11873_new_n1676
* NET  1046 = abc_11873_new_n1675
* NET  1047 = abc_11873_new_n1674
* NET  1048 = abc_11873_new_n1673
* NET  1049 = abc_11873_new_n1672
* NET  1050 = abc_11873_new_n1670
* NET  1051 = abc_11873_new_n1669
* NET  1052 = abc_11873_new_n1668
* NET  1053 = abc_11873_new_n1667
* NET  1054 = abc_11873_new_n1666
* NET  1055 = abc_11873_new_n1665
* NET  1056 = abc_11873_new_n1664
* NET  1057 = abc_11873_new_n1663
* NET  1058 = abc_11873_new_n1662
* NET  1059 = abc_11873_new_n1661
* NET  1060 = abc_11873_new_n1660
* NET  1061 = abc_11873_new_n1658
* NET  1062 = abc_11873_new_n1657
* NET  1063 = abc_11873_new_n1656
* NET  1064 = abc_11873_new_n1655
* NET  1065 = abc_11873_new_n1654
* NET  1066 = abc_11873_new_n1653
* NET  1067 = abc_11873_new_n1652
* NET  1068 = abc_11873_new_n1651
* NET  1069 = abc_11873_new_n1649
* NET  1070 = abc_11873_new_n1648
* NET  1071 = abc_11873_new_n1647
* NET  1072 = abc_11873_new_n1646
* NET  1073 = abc_11873_new_n1645
* NET  1074 = abc_11873_new_n1644
* NET  1075 = abc_11873_new_n1643
* NET  1076 = abc_11873_new_n1642
* NET  1077 = abc_11873_new_n1640
* NET  1078 = abc_11873_new_n1639
* NET  1079 = abc_11873_new_n1638
* NET  1080 = abc_11873_new_n1637
* NET  1081 = abc_11873_new_n1636
* NET  1082 = abc_11873_new_n1635
* NET  1083 = abc_11873_new_n1634
* NET  1084 = abc_11873_new_n1633
* NET  1085 = abc_11873_new_n1632
* NET  1086 = abc_11873_new_n1630
* NET  1087 = abc_11873_new_n1629
* NET  1088 = abc_11873_new_n1628
* NET  1089 = abc_11873_new_n1627
* NET  1090 = abc_11873_new_n1626
* NET  1091 = abc_11873_new_n1625
* NET  1092 = abc_11873_new_n1624
* NET  1093 = abc_11873_new_n1623
* NET  1094 = abc_11873_new_n1622
* NET  1095 = abc_11873_new_n1620
* NET  1096 = abc_11873_new_n1619
* NET  1097 = abc_11873_new_n1618
* NET  1098 = abc_11873_new_n1617
* NET  1099 = abc_11873_new_n1616
* NET  1100 = abc_11873_new_n1615
* NET  1101 = abc_11873_new_n1614
* NET  1102 = abc_11873_new_n1613
* NET  1103 = abc_11873_new_n1611
* NET  1104 = abc_11873_new_n1610
* NET  1105 = abc_11873_new_n1609
* NET  1106 = abc_11873_new_n1608
* NET  1107 = abc_11873_new_n1607
* NET  1108 = abc_11873_new_n1606
* NET  1109 = abc_11873_new_n1605
* NET  1110 = abc_11873_new_n1604
* NET  1111 = abc_11873_new_n1603
* NET  1112 = abc_11873_new_n1602
* NET  1113 = abc_11873_new_n1601
* NET  1114 = abc_11873_new_n1599
* NET  1115 = abc_11873_new_n1598
* NET  1116 = abc_11873_new_n1597
* NET  1117 = abc_11873_new_n1596
* NET  1118 = abc_11873_new_n1595
* NET  1119 = abc_11873_new_n1594
* NET  1120 = abc_11873_new_n1593
* NET  1121 = abc_11873_new_n1592
* NET  1122 = abc_11873_new_n1590
* NET  1123 = abc_11873_new_n1589
* NET  1124 = abc_11873_new_n1588
* NET  1125 = abc_11873_new_n1587
* NET  1126 = abc_11873_new_n1586
* NET  1127 = abc_11873_new_n1585
* NET  1128 = abc_11873_new_n1584
* NET  1129 = abc_11873_new_n1583
* NET  1130 = abc_11873_new_n1582
* NET  1131 = abc_11873_new_n1581
* NET  1132 = abc_11873_new_n1580
* NET  1133 = abc_11873_new_n1579
* NET  1134 = abc_11873_new_n1578
* NET  1135 = abc_11873_new_n1577
* NET  1136 = abc_11873_new_n1576
* NET  1137 = abc_11873_new_n1575
* NET  1138 = abc_11873_new_n1574
* NET  1139 = abc_11873_new_n1573
* NET  1140 = abc_11873_new_n1572
* NET  1141 = abc_11873_new_n1571
* NET  1142 = abc_11873_new_n1570
* NET  1143 = abc_11873_new_n1569
* NET  1144 = abc_11873_new_n1568
* NET  1145 = abc_11873_new_n1551
* NET  1146 = abc_11873_new_n1550
* NET  1147 = abc_11873_new_n1549
* NET  1148 = abc_11873_new_n1548
* NET  1149 = abc_11873_new_n1547
* NET  1150 = abc_11873_new_n1546
* NET  1151 = abc_11873_new_n1545
* NET  1152 = abc_11873_new_n1544
* NET  1153 = abc_11873_new_n1543
* NET  1154 = abc_11873_new_n1542
* NET  1155 = abc_11873_new_n1541
* NET  1156 = abc_11873_new_n1540
* NET  1157 = abc_11873_new_n1539
* NET  1158 = abc_11873_new_n1538
* NET  1159 = abc_11873_new_n1537
* NET  1160 = abc_11873_new_n1536
* NET  1161 = abc_11873_new_n1535
* NET  1162 = abc_11873_new_n1534
* NET  1163 = abc_11873_new_n1533
* NET  1164 = abc_11873_new_n1532
* NET  1165 = abc_11873_new_n1531
* NET  1166 = abc_11873_new_n1530
* NET  1167 = abc_11873_new_n1529
* NET  1168 = abc_11873_new_n1528
* NET  1169 = abc_11873_new_n1527
* NET  1170 = abc_11873_new_n1526
* NET  1171 = abc_11873_new_n1525
* NET  1172 = abc_11873_new_n1524
* NET  1173 = abc_11873_new_n1523
* NET  1174 = abc_11873_new_n1522
* NET  1175 = abc_11873_new_n1521
* NET  1176 = abc_11873_new_n1520
* NET  1177 = abc_11873_new_n1519
* NET  1178 = abc_11873_new_n1518
* NET  1179 = abc_11873_new_n1517
* NET  1180 = abc_11873_new_n1516
* NET  1181 = abc_11873_new_n1515
* NET  1182 = abc_11873_new_n1514
* NET  1183 = abc_11873_new_n1513
* NET  1184 = abc_11873_new_n1512
* NET  1185 = abc_11873_new_n1511
* NET  1186 = abc_11873_new_n1510
* NET  1187 = abc_11873_new_n1509
* NET  1188 = abc_11873_new_n1508
* NET  1189 = abc_11873_new_n1507
* NET  1190 = abc_11873_new_n1506
* NET  1191 = abc_11873_new_n1505
* NET  1192 = abc_11873_new_n1504
* NET  1193 = abc_11873_new_n1503
* NET  1194 = abc_11873_new_n1502
* NET  1195 = abc_11873_new_n1499
* NET  1196 = abc_11873_new_n1498
* NET  1197 = abc_11873_new_n1497
* NET  1198 = abc_11873_new_n1496
* NET  1199 = abc_11873_new_n1495
* NET  1200 = abc_11873_new_n1494
* NET  1201 = abc_11873_new_n1493
* NET  1202 = abc_11873_new_n1492
* NET  1203 = abc_11873_new_n1491
* NET  1204 = abc_11873_new_n1489
* NET  1205 = abc_11873_new_n1488
* NET  1206 = abc_11873_new_n1487
* NET  1207 = abc_11873_new_n1486
* NET  1208 = abc_11873_new_n1485
* NET  1209 = abc_11873_new_n1484
* NET  1210 = abc_11873_new_n1483
* NET  1211 = abc_11873_new_n1482
* NET  1212 = abc_11873_new_n1481
* NET  1213 = abc_11873_new_n1479
* NET  1214 = abc_11873_new_n1478
* NET  1215 = abc_11873_new_n1477
* NET  1216 = abc_11873_new_n1476
* NET  1217 = abc_11873_new_n1475
* NET  1218 = abc_11873_new_n1474
* NET  1219 = abc_11873_new_n1473
* NET  1220 = abc_11873_new_n1471
* NET  1221 = abc_11873_new_n1470
* NET  1222 = abc_11873_new_n1469
* NET  1223 = abc_11873_new_n1468
* NET  1224 = abc_11873_new_n1466
* NET  1225 = abc_11873_new_n1465
* NET  1226 = abc_11873_new_n1464
* NET  1227 = abc_11873_new_n1463
* NET  1228 = abc_11873_new_n1462
* NET  1229 = abc_11873_new_n1461
* NET  1230 = abc_11873_new_n1460
* NET  1231 = abc_11873_new_n1459
* NET  1232 = abc_11873_new_n1457
* NET  1233 = abc_11873_new_n1456
* NET  1234 = abc_11873_new_n1455
* NET  1235 = abc_11873_new_n1454
* NET  1236 = abc_11873_new_n1453
* NET  1237 = abc_11873_new_n1452
* NET  1238 = abc_11873_new_n1451
* NET  1239 = abc_11873_new_n1450
* NET  1240 = abc_11873_new_n1449
* NET  1241 = abc_11873_new_n1448
* NET  1242 = abc_11873_new_n1447
* NET  1243 = abc_11873_new_n1446
* NET  1244 = abc_11873_new_n1436
* NET  1245 = abc_11873_new_n1435
* NET  1246 = abc_11873_new_n1434
* NET  1247 = abc_11873_new_n1432
* NET  1248 = abc_11873_new_n1431
* NET  1249 = abc_11873_new_n1430
* NET  1250 = abc_11873_new_n1429
* NET  1251 = abc_11873_new_n1428
* NET  1252 = abc_11873_new_n1427
* NET  1253 = abc_11873_new_n1426
* NET  1254 = abc_11873_new_n1425
* NET  1255 = abc_11873_new_n1424
* NET  1256 = abc_11873_new_n1423
* NET  1257 = abc_11873_new_n1420
* NET  1258 = abc_11873_new_n1419
* NET  1259 = abc_11873_new_n1418
* NET  1260 = abc_11873_new_n1417
* NET  1261 = abc_11873_new_n1416
* NET  1262 = abc_11873_new_n1414
* NET  1263 = abc_11873_new_n1413
* NET  1264 = abc_11873_new_n1412
* NET  1265 = abc_11873_new_n1411
* NET  1266 = abc_11873_new_n1410
* NET  1267 = abc_11873_new_n1409
* NET  1268 = abc_11873_new_n1407
* NET  1269 = abc_11873_new_n1406
* NET  1270 = abc_11873_new_n1405
* NET  1271 = abc_11873_new_n1404
* NET  1272 = abc_11873_new_n1403
* NET  1273 = abc_11873_new_n1402
* NET  1274 = abc_11873_new_n1401
* NET  1275 = abc_11873_new_n1399
* NET  1276 = abc_11873_new_n1398
* NET  1277 = abc_11873_new_n1397
* NET  1278 = abc_11873_new_n1396
* NET  1279 = abc_11873_new_n1395
* NET  1280 = abc_11873_new_n1394
* NET  1281 = abc_11873_new_n1393
* NET  1282 = abc_11873_new_n1392
* NET  1283 = abc_11873_new_n1391
* NET  1284 = abc_11873_new_n1390
* NET  1285 = abc_11873_new_n1388
* NET  1286 = abc_11873_new_n1387
* NET  1287 = abc_11873_new_n1386
* NET  1288 = abc_11873_new_n1384
* NET  1289 = abc_11873_new_n1383
* NET  1290 = abc_11873_new_n1382
* NET  1291 = abc_11873_new_n1380
* NET  1292 = abc_11873_new_n1378
* NET  1293 = abc_11873_new_n1376
* NET  1294 = abc_11873_new_n1375
* NET  1295 = abc_11873_new_n1374
* NET  1296 = abc_11873_new_n1373
* NET  1297 = abc_11873_new_n1372
* NET  1298 = abc_11873_new_n1369
* NET  1299 = abc_11873_new_n1367
* NET  1300 = abc_11873_new_n1366
* NET  1301 = abc_11873_new_n1365
* NET  1302 = abc_11873_new_n1364
* NET  1303 = abc_11873_new_n1363
* NET  1304 = abc_11873_new_n1362
* NET  1305 = abc_11873_new_n1361
* NET  1306 = abc_11873_new_n1359
* NET  1307 = abc_11873_new_n1358
* NET  1308 = abc_11873_new_n1357
* NET  1309 = abc_11873_new_n1354
* NET  1310 = abc_11873_new_n1353
* NET  1311 = abc_11873_new_n1352
* NET  1312 = abc_11873_new_n1351
* NET  1313 = abc_11873_new_n1350
* NET  1314 = abc_11873_new_n1347
* NET  1315 = abc_11873_new_n1345
* NET  1316 = abc_11873_new_n1344
* NET  1317 = abc_11873_new_n1343
* NET  1318 = abc_11873_new_n1342
* NET  1319 = abc_11873_new_n1341
* NET  1320 = abc_11873_new_n1339
* NET  1321 = abc_11873_new_n1338
* NET  1322 = abc_11873_new_n1337
* NET  1323 = abc_11873_new_n1336
* NET  1324 = abc_11873_new_n1335
* NET  1325 = abc_11873_new_n1334
* NET  1326 = abc_11873_new_n1333
* NET  1327 = abc_11873_new_n1332
* NET  1328 = abc_11873_new_n1331
* NET  1329 = abc_11873_new_n1330
* NET  1330 = abc_11873_new_n1329
* NET  1331 = abc_11873_new_n1328
* NET  1332 = abc_11873_new_n1327
* NET  1333 = abc_11873_new_n1326
* NET  1334 = abc_11873_new_n1325
* NET  1335 = abc_11873_new_n1324
* NET  1336 = abc_11873_new_n1323
* NET  1337 = abc_11873_new_n1322
* NET  1338 = abc_11873_new_n1321
* NET  1339 = abc_11873_new_n1320
* NET  1340 = abc_11873_new_n1319
* NET  1341 = abc_11873_new_n1318
* NET  1342 = abc_11873_new_n1317
* NET  1343 = abc_11873_new_n1316
* NET  1344 = abc_11873_new_n1315
* NET  1345 = abc_11873_new_n1314
* NET  1346 = abc_11873_new_n1313
* NET  1347 = abc_11873_new_n1311
* NET  1348 = abc_11873_new_n1310
* NET  1349 = abc_11873_new_n1308
* NET  1350 = abc_11873_new_n1307
* NET  1351 = abc_11873_new_n1306
* NET  1352 = abc_11873_new_n1305
* NET  1353 = abc_11873_new_n1303
* NET  1354 = abc_11873_new_n1302
* NET  1355 = abc_11873_new_n1300
* NET  1356 = abc_11873_new_n1299
* NET  1357 = abc_11873_new_n1297
* NET  1358 = abc_11873_new_n1296
* NET  1359 = abc_11873_new_n1294
* NET  1360 = abc_11873_new_n1293
* NET  1361 = abc_11873_new_n1292
* NET  1362 = abc_11873_new_n1290
* NET  1363 = abc_11873_new_n1289
* NET  1364 = abc_11873_new_n1287
* NET  1365 = abc_11873_new_n1286
* NET  1366 = abc_11873_new_n1285
* NET  1367 = abc_11873_new_n1283
* NET  1368 = abc_11873_new_n1282
* NET  1369 = abc_11873_new_n1280
* NET  1370 = abc_11873_new_n1279
* NET  1371 = abc_11873_new_n1278
* NET  1372 = abc_11873_new_n1273
* NET  1373 = abc_11873_new_n1264
* NET  1374 = abc_11873_new_n1255
* NET  1375 = abc_11873_new_n1246
* NET  1376 = abc_11873_new_n1244
* NET  1377 = abc_11873_new_n1243
* NET  1378 = abc_11873_new_n1242
* NET  1379 = abc_11873_new_n1241
* NET  1380 = abc_11873_new_n1239
* NET  1381 = abc_11873_new_n1238
* NET  1382 = abc_11873_new_n1237
* NET  1383 = abc_11873_new_n1236
* NET  1384 = abc_11873_new_n1235
* NET  1385 = abc_11873_new_n1233
* NET  1386 = abc_11873_new_n1232
* NET  1387 = abc_11873_new_n1231
* NET  1388 = abc_11873_new_n1230
* NET  1389 = abc_11873_new_n1229
* NET  1390 = abc_11873_new_n1228
* NET  1391 = abc_11873_new_n1227
* NET  1392 = abc_11873_new_n1226
* NET  1393 = abc_11873_new_n1224
* NET  1394 = abc_11873_new_n1222
* NET  1395 = abc_11873_new_n1221
* NET  1396 = abc_11873_new_n1220
* NET  1397 = abc_11873_new_n1219
* NET  1398 = abc_11873_new_n1217
* NET  1399 = abc_11873_new_n1216
* NET  1400 = abc_11873_new_n1215
* NET  1401 = abc_11873_new_n1214
* NET  1402 = abc_11873_new_n1213
* NET  1403 = abc_11873_new_n1211
* NET  1404 = abc_11873_new_n1210
* NET  1405 = abc_11873_new_n1209
* NET  1406 = abc_11873_new_n1208
* NET  1407 = abc_11873_new_n1207
* NET  1408 = abc_11873_new_n1206
* NET  1409 = abc_11873_new_n1205
* NET  1410 = abc_11873_new_n1204
* NET  1411 = abc_11873_new_n1203
* NET  1412 = abc_11873_new_n1201
* NET  1413 = abc_11873_new_n1200
* NET  1414 = abc_11873_new_n1199
* NET  1415 = abc_11873_new_n1198
* NET  1416 = abc_11873_new_n1197
* NET  1417 = abc_11873_new_n1196
* NET  1418 = abc_11873_new_n1195
* NET  1419 = abc_11873_new_n1194
* NET  1420 = abc_11873_new_n1191
* NET  1421 = abc_11873_new_n1190
* NET  1422 = abc_11873_new_n1189
* NET  1423 = abc_11873_new_n1188
* NET  1424 = abc_11873_new_n1187
* NET  1425 = abc_11873_new_n1185
* NET  1426 = abc_11873_new_n1184
* NET  1427 = abc_11873_new_n1183
* NET  1428 = abc_11873_new_n1182
* NET  1429 = abc_11873_new_n1181
* NET  1430 = abc_11873_new_n1179
* NET  1431 = abc_11873_new_n1178
* NET  1432 = abc_11873_new_n1177
* NET  1433 = abc_11873_new_n1176
* NET  1434 = abc_11873_new_n1175
* NET  1435 = abc_11873_new_n1173
* NET  1436 = abc_11873_new_n1172
* NET  1437 = abc_11873_new_n1171
* NET  1438 = abc_11873_new_n1170
* NET  1439 = abc_11873_new_n1169
* NET  1440 = abc_11873_new_n1167
* NET  1441 = abc_11873_new_n1166
* NET  1442 = abc_11873_new_n1165
* NET  1443 = abc_11873_new_n1164
* NET  1444 = abc_11873_new_n1163
* NET  1445 = abc_11873_new_n1161
* NET  1446 = abc_11873_new_n1160
* NET  1447 = abc_11873_new_n1159
* NET  1448 = abc_11873_new_n1158
* NET  1449 = abc_11873_new_n1157
* NET  1450 = abc_11873_new_n1155
* NET  1451 = abc_11873_new_n1154
* NET  1452 = abc_11873_new_n1153
* NET  1453 = abc_11873_new_n1152
* NET  1454 = abc_11873_new_n1151
* NET  1455 = abc_11873_new_n1149
* NET  1456 = abc_11873_new_n1148
* NET  1457 = abc_11873_new_n1147
* NET  1458 = abc_11873_new_n1146
* NET  1459 = abc_11873_new_n1145
* NET  1460 = abc_11873_new_n1144
* NET  1461 = abc_11873_new_n1142
* NET  1462 = abc_11873_new_n1141
* NET  1463 = abc_11873_new_n1140
* NET  1464 = abc_11873_new_n1139
* NET  1465 = abc_11873_new_n1138
* NET  1466 = abc_11873_new_n1137
* NET  1467 = abc_11873_new_n1136
* NET  1468 = abc_11873_new_n1134
* NET  1469 = abc_11873_new_n1133
* NET  1470 = abc_11873_new_n1132
* NET  1471 = abc_11873_new_n1131
* NET  1472 = abc_11873_new_n1130
* NET  1473 = abc_11873_new_n1129
* NET  1474 = abc_11873_new_n1128
* NET  1475 = abc_11873_new_n1126
* NET  1476 = abc_11873_new_n1125
* NET  1477 = abc_11873_new_n1124
* NET  1478 = abc_11873_new_n1123
* NET  1479 = abc_11873_new_n1122
* NET  1480 = abc_11873_new_n1121
* NET  1481 = abc_11873_new_n1120
* NET  1482 = abc_11873_new_n1119
* NET  1483 = abc_11873_new_n1117
* NET  1484 = abc_11873_new_n1116
* NET  1485 = abc_11873_new_n1115
* NET  1486 = abc_11873_new_n1114
* NET  1487 = abc_11873_new_n1113
* NET  1488 = abc_11873_new_n1112
* NET  1489 = abc_11873_new_n1111
* NET  1490 = abc_11873_new_n1109
* NET  1491 = abc_11873_new_n1108
* NET  1492 = abc_11873_new_n1107
* NET  1493 = abc_11873_new_n1106
* NET  1494 = abc_11873_new_n1105
* NET  1495 = abc_11873_new_n1104
* NET  1496 = abc_11873_new_n1103
* NET  1497 = abc_11873_new_n1101
* NET  1498 = abc_11873_new_n1100
* NET  1499 = abc_11873_new_n1099
* NET  1500 = abc_11873_new_n1098
* NET  1501 = abc_11873_new_n1097
* NET  1502 = abc_11873_new_n1096
* NET  1503 = abc_11873_new_n1095
* NET  1504 = abc_11873_new_n1093
* NET  1505 = abc_11873_new_n1092
* NET  1506 = abc_11873_new_n1091
* NET  1507 = abc_11873_new_n1090
* NET  1508 = abc_11873_new_n1089
* NET  1509 = abc_11873_new_n1088
* NET  1510 = abc_11873_new_n1087
* NET  1511 = abc_11873_new_n1085
* NET  1512 = abc_11873_new_n1084
* NET  1513 = abc_11873_new_n1083
* NET  1514 = abc_11873_new_n1082
* NET  1515 = abc_11873_new_n1081
* NET  1516 = abc_11873_new_n1080
* NET  1517 = abc_11873_new_n1079
* NET  1518 = abc_11873_new_n1078
* NET  1519 = abc_11873_new_n1077
* NET  1520 = abc_11873_new_n1076
* NET  1521 = abc_11873_new_n1075
* NET  1522 = abc_11873_new_n1074
* NET  1523 = abc_11873_new_n1073
* NET  1524 = abc_11873_new_n1072
* NET  1525 = abc_11873_new_n1071
* NET  1526 = abc_11873_new_n1070
* NET  1527 = abc_11873_new_n1069
* NET  1528 = abc_11873_new_n1068
* NET  1529 = abc_11873_new_n1067
* NET  1530 = abc_11873_new_n1066
* NET  1531 = abc_11873_new_n1065
* NET  1532 = abc_11873_new_n1064
* NET  1533 = abc_11873_new_n1063
* NET  1534 = abc_11873_new_n1062
* NET  1535 = abc_11873_new_n1061
* NET  1536 = abc_11873_new_n1060
* NET  1537 = abc_11873_new_n1059
* NET  1538 = abc_11873_new_n1058
* NET  1539 = abc_11873_new_n1057
* NET  1540 = abc_11873_new_n1056
* NET  1541 = abc_11873_new_n1055
* NET  1542 = abc_11873_new_n1054
* NET  1543 = abc_11873_new_n1053
* NET  1544 = abc_11873_new_n1052
* NET  1545 = abc_11873_new_n1050
* NET  1546 = abc_11873_new_n1049
* NET  1547 = abc_11873_new_n1048
* NET  1548 = abc_11873_new_n1047
* NET  1549 = abc_11873_new_n1046
* NET  1550 = abc_11873_new_n1045
* NET  1551 = abc_11873_new_n1044
* NET  1552 = abc_11873_new_n1043
* NET  1553 = abc_11873_new_n1042
* NET  1554 = abc_11873_new_n1041
* NET  1555 = abc_11873_new_n1040
* NET  1556 = abc_11873_new_n1038
* NET  1557 = abc_11873_new_n1037
* NET  1558 = abc_11873_new_n1036
* NET  1559 = abc_11873_new_n1035
* NET  1560 = abc_11873_new_n1034
* NET  1561 = abc_11873_new_n1033
* NET  1562 = abc_11873_new_n1032
* NET  1563 = abc_11873_new_n1031
* NET  1564 = abc_11873_new_n1030
* NET  1565 = abc_11873_new_n1029
* NET  1566 = abc_11873_new_n1028
* NET  1567 = abc_11873_new_n1026
* NET  1568 = abc_11873_new_n1025
* NET  1569 = abc_11873_new_n1024
* NET  1570 = abc_11873_new_n1023
* NET  1571 = abc_11873_new_n1022
* NET  1572 = abc_11873_new_n1021
* NET  1573 = abc_11873_new_n1020
* NET  1574 = abc_11873_new_n1019
* NET  1575 = abc_11873_new_n1018
* NET  1576 = abc_11873_new_n1017
* NET  1577 = abc_11873_new_n1016
* NET  1578 = abc_11873_new_n1015
* NET  1579 = abc_11873_new_n1013
* NET  1580 = abc_11873_new_n1012
* NET  1581 = abc_11873_new_n1011
* NET  1582 = abc_11873_new_n1010
* NET  1583 = abc_11873_new_n1009
* NET  1584 = abc_11873_new_n1008
* NET  1585 = abc_11873_new_n1007
* NET  1586 = abc_11873_new_n1006
* NET  1587 = abc_11873_new_n1005
* NET  1588 = abc_11873_new_n1004
* NET  1589 = abc_11873_new_n1003
* NET  1590 = abc_11873_new_n1001
* NET  1591 = abc_11873_new_n1000
* NET  1592 = abc_11873_flatten_MOS6502_0_adj_bcd_0_0
* NET  1593 = abc_11873_auto_rtlil_cc_2560_MuxGate_11872
* NET  1594 = abc_11873_auto_rtlil_cc_2560_MuxGate_11870
* NET  1595 = abc_11873_auto_rtlil_cc_2560_MuxGate_11868
* NET  1596 = abc_11873_auto_rtlil_cc_2560_MuxGate_11866
* NET  1597 = abc_11873_auto_rtlil_cc_2560_MuxGate_11864
* NET  1598 = abc_11873_auto_rtlil_cc_2560_MuxGate_11862
* NET  1599 = abc_11873_auto_rtlil_cc_2560_MuxGate_11860
* NET  1600 = abc_11873_auto_rtlil_cc_2560_MuxGate_11858
* NET  1601 = abc_11873_auto_rtlil_cc_2560_MuxGate_11856
* NET  1602 = abc_11873_auto_rtlil_cc_2560_MuxGate_11854
* NET  1603 = abc_11873_auto_rtlil_cc_2560_MuxGate_11852
* NET  1604 = abc_11873_auto_rtlil_cc_2560_MuxGate_11850
* NET  1605 = abc_11873_auto_rtlil_cc_2560_MuxGate_11848
* NET  1606 = abc_11873_auto_rtlil_cc_2560_MuxGate_11846
* NET  1607 = abc_11873_auto_rtlil_cc_2560_MuxGate_11844
* NET  1608 = abc_11873_auto_rtlil_cc_2560_MuxGate_11842
* NET  1609 = abc_11873_auto_rtlil_cc_2560_MuxGate_11840
* NET  1610 = abc_11873_auto_rtlil_cc_2560_MuxGate_11838
* NET  1611 = abc_11873_auto_rtlil_cc_2560_MuxGate_11836
* NET  1612 = abc_11873_auto_rtlil_cc_2560_MuxGate_11834
* NET  1613 = abc_11873_auto_rtlil_cc_2560_MuxGate_11832
* NET  1614 = abc_11873_auto_rtlil_cc_2560_MuxGate_11830
* NET  1615 = abc_11873_auto_rtlil_cc_2560_MuxGate_11828
* NET  1616 = abc_11873_auto_rtlil_cc_2560_MuxGate_11826
* NET  1617 = abc_11873_auto_rtlil_cc_2560_MuxGate_11824
* NET  1618 = abc_11873_auto_rtlil_cc_2560_MuxGate_11822
* NET  1619 = abc_11873_auto_rtlil_cc_2560_MuxGate_11820
* NET  1620 = abc_11873_auto_rtlil_cc_2560_MuxGate_11818
* NET  1621 = abc_11873_auto_rtlil_cc_2560_MuxGate_11816
* NET  1622 = abc_11873_auto_rtlil_cc_2560_MuxGate_11814
* NET  1623 = abc_11873_auto_rtlil_cc_2560_MuxGate_11812
* NET  1624 = abc_11873_auto_rtlil_cc_2560_MuxGate_11810
* NET  1625 = abc_11873_auto_rtlil_cc_2560_MuxGate_11808
* NET  1626 = abc_11873_auto_rtlil_cc_2560_MuxGate_11806
* NET  1627 = abc_11873_auto_rtlil_cc_2560_MuxGate_11804
* NET  1628 = abc_11873_auto_rtlil_cc_2560_MuxGate_11802
* NET  1629 = abc_11873_auto_rtlil_cc_2560_MuxGate_11800
* NET  1630 = abc_11873_auto_rtlil_cc_2560_MuxGate_11798
* NET  1631 = abc_11873_auto_rtlil_cc_2560_MuxGate_11796
* NET  1632 = abc_11873_auto_rtlil_cc_2560_MuxGate_11794
* NET  1633 = abc_11873_auto_rtlil_cc_2560_MuxGate_11792
* NET  1634 = abc_11873_auto_rtlil_cc_2560_MuxGate_11790
* NET  1635 = abc_11873_auto_rtlil_cc_2560_MuxGate_11788
* NET  1636 = abc_11873_auto_rtlil_cc_2560_MuxGate_11786
* NET  1637 = abc_11873_auto_rtlil_cc_2560_MuxGate_11784
* NET  1638 = abc_11873_auto_rtlil_cc_2560_MuxGate_11782
* NET  1639 = abc_11873_auto_rtlil_cc_2560_MuxGate_11780
* NET  1640 = abc_11873_auto_rtlil_cc_2560_MuxGate_11778
* NET  1641 = abc_11873_auto_rtlil_cc_2560_MuxGate_11776
* NET  1642 = abc_11873_auto_rtlil_cc_2560_MuxGate_11774
* NET  1643 = abc_11873_auto_rtlil_cc_2560_MuxGate_11770
* NET  1644 = abc_11873_auto_rtlil_cc_2560_MuxGate_11768
* NET  1645 = abc_11873_auto_rtlil_cc_2560_MuxGate_11766
* NET  1646 = abc_11873_auto_rtlil_cc_2560_MuxGate_11764
* NET  1647 = abc_11873_auto_rtlil_cc_2560_MuxGate_11762
* NET  1648 = abc_11873_auto_rtlil_cc_2560_MuxGate_11760
* NET  1649 = abc_11873_auto_rtlil_cc_2560_MuxGate_11758
* NET  1650 = abc_11873_auto_rtlil_cc_2560_MuxGate_11756
* NET  1651 = abc_11873_auto_rtlil_cc_2560_MuxGate_11754
* NET  1652 = abc_11873_auto_rtlil_cc_2560_MuxGate_11752
* NET  1653 = abc_11873_auto_rtlil_cc_2560_MuxGate_11748
* NET  1654 = abc_11873_auto_rtlil_cc_2560_MuxGate_11746
* NET  1655 = abc_11873_auto_rtlil_cc_2560_MuxGate_11742
* NET  1656 = abc_11873_auto_rtlil_cc_2560_MuxGate_11740
* NET  1657 = abc_11873_auto_rtlil_cc_2560_MuxGate_11738
* NET  1658 = abc_11873_auto_rtlil_cc_2560_MuxGate_11736
* NET  1659 = abc_11873_auto_rtlil_cc_2560_MuxGate_11734
* NET  1660 = abc_11873_auto_rtlil_cc_2560_MuxGate_11732
* NET  1661 = abc_11873_auto_rtlil_cc_2560_MuxGate_11730
* NET  1662 = abc_11873_auto_rtlil_cc_2560_MuxGate_11728
* NET  1663 = abc_11873_auto_rtlil_cc_2560_MuxGate_11726
* NET  1664 = abc_11873_auto_rtlil_cc_2560_MuxGate_11724
* NET  1665 = abc_11873_auto_rtlil_cc_2560_MuxGate_11722
* NET  1666 = abc_11873_auto_rtlil_cc_2560_MuxGate_11720
* NET  1667 = abc_11873_auto_rtlil_cc_2560_MuxGate_11716
* NET  1668 = abc_11873_auto_rtlil_cc_2560_MuxGate_11714
* NET  1669 = abc_11873_auto_rtlil_cc_2560_MuxGate_11712
* NET  1670 = abc_11873_auto_rtlil_cc_2560_MuxGate_11710
* NET  1671 = abc_11873_auto_rtlil_cc_2560_MuxGate_11708
* NET  1672 = abc_11873_auto_rtlil_cc_2560_MuxGate_11706
* NET  1673 = abc_11873_auto_rtlil_cc_2560_MuxGate_11704
* NET  1674 = abc_11873_auto_rtlil_cc_2560_MuxGate_11702
* NET  1675 = abc_11873_auto_rtlil_cc_2560_MuxGate_11700
* NET  1676 = abc_11873_auto_rtlil_cc_2560_MuxGate_11698
* NET  1677 = abc_11873_auto_rtlil_cc_2560_MuxGate_11696
* NET  1678 = abc_11873_auto_rtlil_cc_2560_MuxGate_11694
* NET  1679 = abc_11873_auto_rtlil_cc_2560_MuxGate_11692
* NET  1680 = abc_11873_auto_rtlil_cc_2560_MuxGate_11690
* NET  1681 = abc_11873_auto_rtlil_cc_2560_MuxGate_11688
* NET  1682 = abc_11873_auto_rtlil_cc_2560_MuxGate_11686
* NET  1683 = abc_11873_auto_rtlil_cc_2560_MuxGate_11684
* NET  1684 = abc_11873_auto_rtlil_cc_2560_MuxGate_11682
* NET  1685 = abc_11873_auto_rtlil_cc_2560_MuxGate_11680
* NET  1686 = abc_11873_auto_rtlil_cc_2560_MuxGate_11678
* NET  1687 = abc_11873_auto_rtlil_cc_2560_MuxGate_11676
* NET  1688 = abc_11873_auto_rtlil_cc_2560_MuxGate_11672
* NET  1689 = abc_11873_auto_rtlil_cc_2560_MuxGate_11670
* NET  1690 = abc_11873_auto_rtlil_cc_2560_MuxGate_11668
* NET  1691 = abc_11873_auto_rtlil_cc_2560_MuxGate_11666
* NET  1692 = abc_11873_auto_rtlil_cc_2560_MuxGate_11664
* NET  1693 = abc_11873_auto_rtlil_cc_2560_MuxGate_11662
* NET  1694 = abc_11873_auto_rtlil_cc_2560_MuxGate_11660
* NET  1695 = abc_11873_auto_rtlil_cc_2560_MuxGate_11658
* NET  1696 = abc_11873_auto_rtlil_cc_2560_MuxGate_11656
* NET  1697 = abc_11873_auto_rtlil_cc_2560_MuxGate_11654
* NET  1698 = abc_11873_auto_rtlil_cc_2560_MuxGate_11652
* NET  1699 = abc_11873_auto_rtlil_cc_2560_MuxGate_11650
* NET  1700 = abc_11873_auto_rtlil_cc_2560_MuxGate_11648
* NET  1701 = abc_11873_auto_rtlil_cc_2560_MuxGate_11646
* NET  1702 = abc_11873_auto_rtlil_cc_2560_MuxGate_11644
* NET  1703 = abc_11873_auto_rtlil_cc_2560_MuxGate_11642
* NET  1704 = abc_11873_auto_rtlil_cc_2560_MuxGate_11640
* NET  1705 = abc_11873_auto_rtlil_cc_2560_MuxGate_11638
* NET  1706 = abc_11873_auto_rtlil_cc_2560_MuxGate_11636
* NET  1707 = abc_11873_auto_rtlil_cc_2560_MuxGate_11634
* NET  1708 = abc_11873_auto_rtlil_cc_2560_MuxGate_11632
* NET  1709 = abc_11873_auto_rtlil_cc_2560_MuxGate_11630
* NET  1710 = abc_11873_auto_rtlil_cc_2560_MuxGate_11628
* NET  1711 = abc_11873_auto_rtlil_cc_2560_MuxGate_11626
* NET  1712 = abc_11873_auto_rtlil_cc_2560_MuxGate_11624
* NET  1713 = abc_11873_auto_rtlil_cc_2560_MuxGate_11622
* NET  1714 = abc_11873_auto_rtlil_cc_2560_MuxGate_11620
* NET  1715 = abc_11873_auto_rtlil_cc_2560_MuxGate_11618
* NET  1716 = abc_11873_auto_rtlil_cc_2560_MuxGate_11616
* NET  1717 = abc_11873_auto_rtlil_cc_2560_MuxGate_11614
* NET  1718 = abc_11873_auto_rtlil_cc_2560_MuxGate_11612
* NET  1719 = abc_11873_auto_rtlil_cc_2560_MuxGate_11610
* NET  1720 = WE
* NET  1721 = RDY
* NET  1722 = NMI
* NET  1723 = MOS6502_write_back
* NET  1724 = MOS6502_store
* NET  1725 = MOS6502_state[5]
* NET  1726 = MOS6502_state[4]
* NET  1727 = MOS6502_state[3]
* NET  1728 = MOS6502_state[2]
* NET  1729 = MOS6502_state[1]
* NET  1730 = MOS6502_state[0]
* NET  1731 = MOS6502_src_reg[1]
* NET  1732 = MOS6502_src_reg[0]
* NET  1733 = MOS6502_shift_right
* NET  1734 = MOS6502_shift
* NET  1735 = MOS6502_sei
* NET  1736 = MOS6502_sed
* NET  1737 = MOS6502_sec
* NET  1738 = MOS6502_rotate
* NET  1739 = MOS6502_res
* NET  1740 = MOS6502_plp
* NET  1741 = MOS6502_php
* NET  1742 = MOS6502_op[3]
* NET  1743 = MOS6502_op[2]
* NET  1744 = MOS6502_op[1]
* NET  1745 = MOS6502_op[0]
* NET  1746 = MOS6502_load_reg
* NET  1747 = MOS6502_load_only
* NET  1748 = MOS6502_index_y
* NET  1749 = MOS6502_inc
* NET  1750 = MOS6502_dst_reg[1]
* NET  1751 = MOS6502_dst_reg[0]
* NET  1752 = MOS6502_cond_code[2]
* NET  1753 = MOS6502_cond_code[1]
* NET  1754 = MOS6502_cond_code[0]
* NET  1755 = MOS6502_compare
* NET  1756 = MOS6502_clv
* NET  1757 = MOS6502_cli
* NET  1758 = MOS6502_cld
* NET  1759 = MOS6502_clc
* NET  1760 = MOS6502_bit_ins
* NET  1761 = MOS6502_backwards
* NET  1762 = MOS6502_adj_bcd
* NET  1763 = MOS6502_adc_sbc
* NET  1764 = MOS6502_adc_bcd
* NET  1765 = MOS6502_Z
* NET  1766 = MOS6502_V
* NET  1767 = MOS6502_PC[9]
* NET  1768 = MOS6502_PC[8]
* NET  1769 = MOS6502_PC[7]
* NET  1770 = MOS6502_PC[6]
* NET  1771 = MOS6502_PC[5]
* NET  1772 = MOS6502_PC[4]
* NET  1773 = MOS6502_PC[3]
* NET  1774 = MOS6502_PC[2]
* NET  1775 = MOS6502_PC[15]
* NET  1776 = MOS6502_PC[14]
* NET  1777 = MOS6502_PC[13]
* NET  1778 = MOS6502_PC[12]
* NET  1779 = MOS6502_PC[11]
* NET  1780 = MOS6502_PC[10]
* NET  1781 = MOS6502_PC[1]
* NET  1782 = MOS6502_PC[0]
* NET  1783 = MOS6502_NMI_edge
* NET  1784 = MOS6502_NMI_1
* NET  1785 = MOS6502_N
* NET  1786 = MOS6502_IRHOLD_valid
* NET  1787 = MOS6502_IRHOLD[7]
* NET  1788 = MOS6502_IRHOLD[6]
* NET  1789 = MOS6502_IRHOLD[5]
* NET  1790 = MOS6502_IRHOLD[4]
* NET  1791 = MOS6502_IRHOLD[3]
* NET  1792 = MOS6502_IRHOLD[2]
* NET  1793 = MOS6502_IRHOLD[1]
* NET  1794 = MOS6502_IRHOLD[0]
* NET  1795 = MOS6502_I
* NET  1796 = MOS6502_DIMUX[7]
* NET  1797 = MOS6502_DIMUX[6]
* NET  1798 = MOS6502_DIMUX[5]
* NET  1799 = MOS6502_DIMUX[4]
* NET  1800 = MOS6502_DIMUX[3]
* NET  1801 = MOS6502_DIMUX[2]
* NET  1802 = MOS6502_DIMUX[1]
* NET  1803 = MOS6502_DIMUX[0]
* NET  1804 = MOS6502_DIHOLD[7]
* NET  1805 = MOS6502_DIHOLD[6]
* NET  1806 = MOS6502_DIHOLD[5]
* NET  1807 = MOS6502_DIHOLD[4]
* NET  1808 = MOS6502_DIHOLD[3]
* NET  1809 = MOS6502_DIHOLD[2]
* NET  1810 = MOS6502_DIHOLD[1]
* NET  1811 = MOS6502_DIHOLD[0]
* NET  1812 = MOS6502_D
* NET  1813 = MOS6502_C
* NET  1814 = MOS6502_AXYS_3_7
* NET  1815 = MOS6502_AXYS_3_6
* NET  1816 = MOS6502_AXYS_3_5
* NET  1817 = MOS6502_AXYS_3_4
* NET  1818 = MOS6502_AXYS_3_3
* NET  1819 = MOS6502_AXYS_3_2
* NET  1820 = MOS6502_AXYS_3_1
* NET  1821 = MOS6502_AXYS_3_0
* NET  1822 = MOS6502_AXYS_2_7
* NET  1823 = MOS6502_AXYS_2_6
* NET  1824 = MOS6502_AXYS_2_5
* NET  1825 = MOS6502_AXYS_2_4
* NET  1826 = MOS6502_AXYS_2_3
* NET  1827 = MOS6502_AXYS_2_2
* NET  1828 = MOS6502_AXYS_2_1
* NET  1829 = MOS6502_AXYS_2_0
* NET  1830 = MOS6502_AXYS_1_7
* NET  1831 = MOS6502_AXYS_1_6
* NET  1832 = MOS6502_AXYS_1_5
* NET  1833 = MOS6502_AXYS_1_4
* NET  1834 = MOS6502_AXYS_1_3
* NET  1835 = MOS6502_AXYS_1_2
* NET  1836 = MOS6502_AXYS_1_1
* NET  1837 = MOS6502_AXYS_1_0
* NET  1838 = MOS6502_AXYS_0_7
* NET  1839 = MOS6502_AXYS_0_6
* NET  1840 = MOS6502_AXYS_0_5
* NET  1841 = MOS6502_AXYS_0_4
* NET  1842 = MOS6502_AXYS_0_3
* NET  1843 = MOS6502_AXYS_0_2
* NET  1844 = MOS6502_AXYS_0_1
* NET  1845 = MOS6502_AXYS_0_0
* NET  1846 = MOS6502_ALU_OUT[7]
* NET  1847 = MOS6502_ALU_OUT[6]
* NET  1848 = MOS6502_ALU_OUT[5]
* NET  1849 = MOS6502_ALU_OUT[4]
* NET  1850 = MOS6502_ALU_OUT[3]
* NET  1851 = MOS6502_ALU_OUT[2]
* NET  1852 = MOS6502_ALU_OUT[1]
* NET  1853 = MOS6502_ALU_OUT[0]
* NET  1854 = MOS6502_ALU_HC
* NET  1855 = MOS6502_ALU_CO
* NET  1856 = MOS6502_ALU_BI7
* NET  1857 = MOS6502_ALU_AI7
* NET  1858 = MOS6502_ABL[7]
* NET  1859 = MOS6502_ABL[6]
* NET  1860 = MOS6502_ABL[5]
* NET  1861 = MOS6502_ABL[4]
* NET  1862 = MOS6502_ABL[3]
* NET  1863 = MOS6502_ABL[2]
* NET  1864 = MOS6502_ABL[1]
* NET  1865 = MOS6502_ABL[0]
* NET  1866 = MOS6502_ABH[7]
* NET  1867 = MOS6502_ABH[6]
* NET  1868 = MOS6502_ABH[5]
* NET  1869 = MOS6502_ABH[4]
* NET  1870 = MOS6502_ABH[3]
* NET  1871 = MOS6502_ABH[2]
* NET  1872 = MOS6502_ABH[1]
* NET  1873 = MOS6502_ABH[0]
* NET  1874 = IRQ
* NET  1875 = DO[7]
* NET  1876 = DO[6]
* NET  1877 = DO[5]
* NET  1878 = DO[4]
* NET  1879 = DO[3]
* NET  1880 = DO[2]
* NET  1881 = DO[1]
* NET  1882 = DO[0]
* NET  1883 = DI[7]
* NET  1884 = DI[6]
* NET  1885 = DI[5]
* NET  1886 = DI[4]
* NET  1887 = DI[3]
* NET  1888 = DI[2]
* NET  1889 = DI[1]
* NET  1890 = DI[0]
* NET  1891 = A[9]
* NET  1892 = A[8]
* NET  1893 = A[7]
* NET  1894 = A[6]
* NET  1895 = A[5]
* NET  1896 = A[4]
* NET  1897 = A[3]
* NET  1898 = A[2]
* NET  1899 = A[15]
* NET  1900 = A[14]
* NET  1901 = A[13]
* NET  1902 = A[12]
* NET  1903 = A[11]
* NET  1904 = A[10]
* NET  1905 = A[1]
* NET  1906 = A[0]

xsubckt_1742_mx2_x2 0 1597 1 656 677 1848 mx2_x2
xsubckt_1741_mx2_x2 0 1598 1 656 671 1849 mx2_x2
xsubckt_1539_a3_x2 1 867 0 932 937 1798 a3_x2
xsubckt_1461_oa22_x2 0 944 1 1550 956 946 oa22_x2
xsubckt_1450_a3_x2 1 955 0 325 360 377 a3_x2
xsubckt_1285_a3_x2 1 1106 0 1107 1115 1124 a3_x2
xsubckt_495_ao22_x2 0 183 1 527 532 550 ao22_x2
xsubckt_465_mx2_x2 0 212 1 1753 213 214 mx2_x2
xsubckt_464_mx2_x2 0 213 1 1752 1785 1813 mx2_x2
xsubckt_463_mx2_x2 0 214 1 1752 1766 1765 mx2_x2
xsubckt_458_o2_x2 0 219 1 320 466 o2_x2
xsubckt_118_mx2_x2 0 557 1 656 599 600 mx2_x2
xsubckt_653_oa22_x2 0 31 1 44 343 639 oa22_x2
xsubckt_663_o2_x2 0 22 1 51 618 o2_x2
xsubckt_821_nand3_x0 1 0 1460 1518 1526 1768 nand3_x0
xsubckt_962_nand2_x0 1 0 1366 438 1759 nand2_x0
xsubckt_1858_sff1_x4 1 9 0 1626 1871 sff1_x4
xsubckt_1819_sff1_x4 1 9 0 1656 1751 sff1_x4
xsubckt_1770_sff1_x4 1 9 0 3 1725 sff1_x4
xsubckt_1744_mx2_x2 0 1595 1 656 678 1846 mx2_x2
xsubckt_1743_mx2_x2 0 1596 1 656 676 1847 mx2_x2
xsubckt_1569_a3_x2 1 837 0 481 554 1772 a3_x2
xsubckt_1343_a2_x2 0 1054 1 1055 1059 a2_x2
xsubckt_1299_nand3_x0 1 0 1094 545 550 1861 nand3_x0
xsubckt_604_nand2_x0 1 0 79 358 450 nand2_x0
xsubckt_388_nand3_x0 1 0 288 551 588 1727 nand3_x0
xsubckt_337_nand4_x0 1 0 339 467 476 490 554 nand4_x0
xsubckt_995_nand4_x0 1 0 1341 412 517 520 533 nand4_x0
xsubckt_1748_mx2_x2 0 1593 1 656 944 1857 mx2_x2
xsubckt_1667_a2_x2 0 739 1 740 744 a2_x2
xsubckt_1637_a2_x2 0 769 1 771 911 a2_x2
xsubckt_1449_o4_x2 0 956 1 958 959 1172 76 o4_x2
xsubckt_1358_mx2_x2 0 1611 1 656 1041 1767 mx2_x2
xsubckt_1330_oa22_x2 0 1066 1 1846 1135 1067 oa22_x2
xsubckt_727_nand4_x0 1 0 1545 1546 1547 1548 1549 nand4_x0
xsubckt_1766_sff1_x4 1 9 0 7 1729 sff1_x4
xsubckt_1326_nxr2_x1 1069 1 0 1071 1078 nxr2_x1
xsubckt_914_nxr2_x1 1382 1 0 1392 643 nxr2_x1
xsubckt_1672_nand3_x0 1 0 734 932 937 1803 nand3_x0
xsubckt_547_nand4_x0 1 0 132 275 467 1726 587 nand4_x0
xsubckt_1545_nand2_x0 1 0 861 864 911 nand2_x0
xsubckt_582_a4_x2 0 98 1 202 204 225 227 a4_x2
xsubckt_542_a4_x2 0 136 1 137 142 206 228 a4_x2
xsubckt_415_a3_x2 1 261 0 262 298 301 a3_x2
xsubckt_367_nand4_x0 1 0 309 476 490 586 1725 nand4_x0
xsubckt_347_a4_x2 0 329 1 330 333 335 339 a4_x2
xsubckt_281_nand3_x0 1 0 395 467 481 493 nand3_x0
xsubckt_710_nand4_x0 1 0 1561 1563 1564 1565 1566 nand4_x0
xsubckt_988_nand3_x0 1 0 1347 256 404 533 nand3_x0
xsubckt_592_a4_x2 0 89 1 159 160 192 193 a4_x2
xsubckt_445_a3_x2 1 232 0 233 516 520 a3_x2
xsubckt_435_a3_x2 1 242 0 275 586 1725 a3_x2
xsubckt_191_a3_x2 1 485 0 552 590 1729 a3_x2
xsubckt_671_nand3_x0 1 0 15 57 64 1834 nand3_x0
xsubckt_826_a4_x2 0 1455 1 1456 1457 1459 1536 a4_x2
xsubckt_553_a2_x2 0 126 1 127 128 a2_x2
xsubckt_358_a2_x2 0 318 1 319 324 a2_x2
xsubckt_729_a3_x2 1 1544 0 78 85 425 a3_x2
xsubckt_896_oa22_x2 0 1397 1 1406 1401 1402 oa22_x2
xsubckt_1134_nand3_x0 1 0 1232 1233 1235 1236 nand3_x0
xsubckt_1269_oa22_x2 0 1121 1 1131 371 632 oa22_x2
xsubckt_1275_nand2_x0 1 0 1115 1117 1121 nand2_x0
xsubckt_1665_nand2_x0 1 0 741 742 911 nand2_x0
xsubckt_1575_nand2_x0 1 0 831 832 838 nand2_x0
xsubckt_1302_ao22_x2 0 1091 1 646 1136 1093 ao22_x2
xsubckt_573_a2_x2 0 106 1 107 108 a2_x2
xsubckt_368_a2_x2 0 308 1 310 467 a2_x2
xsubckt_881_nand3_x0 1 0 1410 1854 1764 1762 nand3_x0
xsubckt_971_nand3_x0 1 0 1359 1360 1365 412 nand3_x0
xsubckt_994_a3_x2 1 1342 0 517 520 533 a3_x2
xsubckt_1044_nand3_x0 1 0 1299 1300 1301 251 nand3_x0
xsubckt_1210_a4_x2 0 1163 1 1164 1165 1167 1178 a4_x2
xsubckt_1485_nand2_x0 1 0 920 922 977 nand2_x0
xsubckt_397_nand4_x0 1 0 279 551 554 588 1727 nand4_x0
xsubckt_184_nand2_x0 1 0 492 1726 587 nand2_x0
xsubckt_242_oa22_x2 0 434 1 543 541 436 oa22_x2
xsubckt_1882_sff1_x4 1 9 0 1602 1853 sff1_x4
xsubckt_1733_ao22_x2 0 1603 1 674 680 902 ao22_x2
xsubckt_122_nor2_x0 1 0 554 1726 1725 nor2_x0
xsubckt_1843_sff1_x4 1 9 0 1640 1785 sff1_x4
xsubckt_1804_sff1_x4 1 9 0 1671 1743 sff1_x4
xsubckt_1622_a3_x2 1 784 0 932 937 1801 a3_x2
xsubckt_634_oa22_x2 0 49 1 281 360 633 oa22_x2
xsubckt_394_nand2_x0 1 0 282 283 284 nand2_x0
xsubckt_306_nand2_x0 1 0 370 372 467 nand2_x0
xsubckt_823_nand3_x0 1 0 1458 1524 369 482 nand3_x0
xsubckt_1046_a2_x2 0 1298 1 438 1734 a2_x2
xsubckt_1878_sff1_x4 1 9 0 1606 1776 sff1_x4
xsubckt_1839_sff1_x4 1 9 0 1644 1787 sff1_x4
xsubckt_1790_sff1_x4 1 9 0 1685 1753 sff1_x4
xsubckt_1751_sff1_x4 1 9 0 1717 1843 sff1_x4
xsubckt_1684_mx3_x2 1 0 722 977 897 759 725 728 mx3_x2
xsubckt_1683_mx3_x2 1 0 723 977 897 758 724 729 mx3_x2
xsubckt_1487_a3_x2 1 918 0 383 554 1761 a3_x2
xsubckt_1403_oa22_x2 0 999 1 1020 1011 1002 oa22_x2
xsubckt_185_oa22_x2 0 491 1 492 494 498 oa22_x2
xsubckt_253_nand3_x0 1 0 423 467 481 495 nand3_x0
xsubckt_290_nand4_x0 1 0 386 476 587 1728 589 nand4_x0
xsubckt_733_nand3_x0 1 0 1540 1542 351 375 nand3_x0
xsubckt_1477_oa22_x2 0 928 1 1524 460 624 oa22_x2
xsubckt_1464_nand3_x0 1 0 941 942 1524 460 nand3_x0
xsubckt_1337_nand2_x0 1 0 1060 1130 1768 nand2_x0
xsubckt_784_nand2_x0 1 0 1492 1493 1494 nand2_x0
xsubckt_1165_mx2_x2 0 1205 1 377 1802 1852 mx2_x2
xsubckt_1166_mx2_x2 0 1204 1 1209 1205 1206 mx2_x2
xsubckt_1167_mx2_x2 0 1639 1 1211 1765 1204 mx2_x2
xsubckt_1786_sff1_x4 1 9 0 1688 1822 sff1_x4
xsubckt_1307_nxr2_x1 1086 1 0 1089 1096 nxr2_x1
xsubckt_215_a4_x2 0 461 1 552 554 1730 591 a4_x2
xsubckt_776_ao22_x2 0 1499 1 1527 1535 1851 ao22_x2
xsubckt_1016_nand3_x0 1 0 1320 1323 1344 1347 nand3_x0
xsubckt_1067_nand2_x0 1 0 1284 438 584 nand2_x0
xsubckt_1457_nand2_x0 1 0 948 950 984 nand2_x0
xsubckt_1293_oa22_x2 0 1099 1 1850 1135 1100 oa22_x2
xsubckt_539_a4_x2 0 139 1 140 141 313 315 a4_x2
xsubckt_156_nand2_x0 1 0 520 522 523 nand2_x0
xsubckt_4_inv_x0 1 0 1783 664 inv_x0
xsubckt_3_inv_x0 1 0 1812 665 inv_x0
xsubckt_2_inv_x0 1 0 1739 666 inv_x0
xsubckt_1_inv_x0 1 0 1786 667 inv_x0
xsubckt_0_inv_x0 1 0 1795 668 inv_x0
xsubckt_1215_oa22_x2 0 1158 1 494 492 361 oa22_x2
xsubckt_493_nand3_x0 1 0 185 367 383 554 nand3_x0
xsubckt_431_a2_x2 0 246 1 247 252 a2_x2
xsubckt_405_nand3_x0 1 0 271 467 489 493 nand3_x0
xsubckt_9_inv_x0 1 0 1737 659 inv_x0
xsubckt_8_inv_x0 1 0 1740 660 inv_x0
xsubckt_7_inv_x0 1 0 1759 661 inv_x0
xsubckt_6_inv_x0 1 0 1723 662 inv_x0
xsubckt_5_inv_x0 1 0 1734 663 inv_x0
xsubckt_189_nand4_x0 1 0 487 490 1726 1730 591 nand4_x0
xsubckt_256_a2_x2 0 420 1 421 546 a2_x2
xsubckt_315_nand3_x0 1 0 361 476 588 1727 nand3_x0
xsubckt_761_nor2_x0 1 0 1512 1513 1516 nor2_x0
xsubckt_832_a3_x2 1 1450 0 1451 1452 1453 a3_x2
xsubckt_862_a3_x2 1 1425 0 1426 1427 1428 a3_x2
xsubckt_1050_nand2_x0 1 0 1296 438 1749 nand2_x0
xsubckt_1322_ao22_x2 0 1073 1 643 1136 1075 ao22_x2
xsubckt_491_a2_x2 0 186 1 187 303 a2_x2
xsubckt_286_nor3_x0 1 0 390 393 396 426 nor3_x0
xsubckt_705_nand3_x0 1 0 1566 57 63 1815 nand3_x0
xsubckt_745_a2_x2 0 1528 1 1529 369 a2_x2
xsubckt_750_oa22_x2 0 1523 1 495 473 310 oa22_x2
xsubckt_882_a3_x2 1 1409 0 649 650 1762 a3_x2
xsubckt_883_nand3_x0 1 0 1408 649 650 1762 nand3_x0
xsubckt_950_a2_x2 0 1372 1 602 1722 a2_x2
xsubckt_1593_oa22_x2 0 813 1 13 956 815 oa22_x2
xsubckt_1499_nor4_x0 1 0 906 911 918 919 84 nor4_x0
xsubckt_399_nand4_x0 1 0 277 278 280 283 284 nand4_x0
xsubckt_742_nand4_x0 1 0 1531 1534 385 453 471 nand4_x0
xsubckt_900_mx2_x2 0 1716 1 1413 1842 1394 mx2_x2
xsubckt_901_mx2_x2 0 1393 1 354 1799 1849 mx2_x2
xsubckt_1554_oa22_x2 0 852 1 1571 956 854 oa22_x2
xsubckt_1397_nand2_x0 1 0 1005 372 1848 nand2_x0
xsubckt_254_mx3_x2 1 0 422 667 1721 595 596 597 mx3_x2
xsubckt_902_mx2_x2 0 1715 1 1413 1841 1393 mx2_x2
xsubckt_1041_a3_x2 1 1302 0 251 516 521 a3_x2
xsubckt_1219_nand2_x0 1 0 1154 1155 334 nand2_x0
xsubckt_1863_sff1_x4 1 9 0 1621 1866 sff1_x4
xsubckt_1824_sff1_x4 1 9 0 1801 1809 sff1_x4
xsubckt_1714_ao22_x2 0 692 1 701 694 693 ao22_x2
xsubckt_1535_mx3_x2 1 0 871 977 880 945 877 874 mx3_x2
xsubckt_1534_mx3_x2 1 0 872 977 879 944 873 878 mx3_x2
xsubckt_1405_mx2_x2 0 1607 1 656 998 1777 mx2_x2
xsubckt_699_nand4_x0 1 0 1571 1574 1575 1576 1577 nand4_x0
xsubckt_966_nand2_x0 1 0 1363 438 1737 nand2_x0
xsubckt_1080_nand2_x0 1 0 1272 1294 1338 nand2_x0
xsubckt_1142_mx3_x2 1 0 1225 377 240 562 1757 648 mx3_x2
xsubckt_1208_a2_x2 0 1165 1 1166 488 a2_x2
xsubckt_1859_sff1_x4 1 9 0 1625 1870 sff1_x4
xsubckt_1697_nand2_x0 1 0 709 741 743 nand2_x0
xsubckt_1669_a3_x2 1 737 0 481 554 1782 a3_x2
xsubckt_1649_a3_x2 1 757 0 481 554 1781 a3_x2
xsubckt_1463_a2_x2 0 942 1 452 549 a2_x2
xsubckt_1462_oa22_x2 0 943 1 1524 460 625 oa22_x2
xsubckt_1423_a2_x2 0 981 1 982 987 a2_x2
xsubckt_382_nand4_x0 1 0 294 402 404 437 539 nand4_x0
xsubckt_131_oa22_x2 0 545 1 668 1874 1783 oa22_x2
xsubckt_814_ao22_x2 0 1466 1 1527 1535 1846 ao22_x2
xsubckt_1076_nand3_x0 1 0 1275 1276 1279 1334 nand3_x0
xsubckt_1225_o4_x2 0 1148 1 1149 1168 1533 346 o4_x2
xsubckt_1265_ao22_x2 0 1124 1 1125 1127 1139 ao22_x2
xsubckt_1771_sff1_x4 1 9 0 1703 1837 sff1_x4
xsubckt_1727_a2_x2 0 679 1 895 907 a2_x2
xsubckt_1717_a2_x2 0 689 1 690 820 a2_x2
xsubckt_1288_a2_x2 0 1103 1 1104 1105 a2_x2
xsubckt_645_nand3_x0 1 0 39 57 64 1836 nand3_x0
xsubckt_689_oa22_x2 0 1580 1 281 360 629 oa22_x2
xsubckt_786_nand2_x0 1 0 1490 1491 1496 nand2_x0
xsubckt_1173_ao22_x2 0 1198 1 1200 1203 377 ao22_x2
xsubckt_1202_nand2_x0 1 0 1171 1189 270 nand2_x0
xsubckt_1767_sff1_x4 1 9 0 6 1728 sff1_x4
xsubckt_1680_nand2_x0 1 0 726 727 728 nand2_x0
xsubckt_1618_ao22_x2 0 788 1 25 957 790 ao22_x2
xsubckt_1331_oa22_x2 0 1065 1 1769 1128 1066 oa22_x2
xsubckt_1286_nand3_x0 1 0 1105 1107 1115 1124 nand3_x0
xsubckt_10_inv_x0 1 0 1763 658 inv_x0
xsubckt_11_inv_x0 1 0 1755 657 inv_x0
xsubckt_12_inv_x0 1 0 1721 656 inv_x0
xsubckt_13_inv_x0 1 0 2 655 inv_x0
xsubckt_14_inv_x0 1 0 1756 654 inv_x0
xsubckt_1022_nand2_x0 1 0 1315 1316 1318 nand2_x0
xsubckt_375_nand3_x0 1 0 301 467 489 495 nand3_x0
xsubckt_15_inv_x0 1 0 1758 653 inv_x0
xsubckt_16_inv_x0 1 0 1853 652 inv_x0
xsubckt_17_inv_x0 1 0 1852 651 inv_x0
xsubckt_18_inv_x0 1 0 1764 650 inv_x0
xsubckt_19_inv_x0 1 0 1854 649 inv_x0
xsubckt_163_a4_x2 0 513 1 516 521 527 532 a4_x2
xsubckt_234_ao22_x2 0 442 1 443 449 556 ao22_x2
xsubckt_757_ao22_x2 0 1516 1 1527 1535 1853 ao22_x2
xsubckt_796_ao22_x2 0 1482 1 1578 1573 1543 ao22_x2
xsubckt_915_nxr2_x1 1381 1 0 1382 1387 nxr2_x1
xsubckt_996_nand2_x0 1 0 1340 1341 514 nand2_x0
xsubckt_1069_nand2_x0 1 0 1282 1283 1326 nand2_x0
xsubckt_1586_nand3_x0 1 0 820 821 826 841 nand3_x0
xsubckt_1526_ao22_x2 0 880 1 1562 957 882 ao22_x2
xsubckt_501_nand2_x0 1 0 177 505 538 nand2_x0
xsubckt_466_nxr2_x1 211 1 0 212 640 nxr2_x1
xsubckt_765_nand3_x0 1 0 1509 1518 1526 1781 nand3_x0
xsubckt_1496_nand3_x0 1 0 909 911 913 914 nand3_x0
xsubckt_142_ao22_x2 0 534 1 1786 1801 546 ao22_x2
xsubckt_134_a2_x2 0 542 1 543 546 a2_x2
xsubckt_124_a2_x2 0 552 1 1728 1727 a2_x2
xsubckt_269_ao22_x2 0 407 1 414 418 420 ao22_x2
xsubckt_284_nor4_x0 1 0 392 393 428 433 440 nor4_x0
xsubckt_672_a4_x2 0 14 1 15 16 17 18 a4_x2
xsubckt_897_nxr2_x1 1396 1 0 1409 1850 nxr2_x1
xsubckt_555_a3_x2 1 124 0 125 140 141 a3_x2
xsubckt_317_nand3_x0 1 0 359 362 467 493 nand3_x0
xsubckt_770_a3_x2 1 1504 0 1505 1508 1509 a3_x2
xsubckt_801_nand2_x0 1 0 1477 1478 1479 nand2_x0
xsubckt_1666_oa22_x2 0 740 1 911 742 906 oa22_x2
xsubckt_1627_oa22_x2 0 779 1 783 785 939 oa22_x2
xsubckt_488_a2_x2 0 189 1 190 195 a2_x2
xsubckt_354_nand4_x0 1 0 322 552 587 590 1729 nand4_x0
xsubckt_707_nand3_x0 1 0 1564 57 64 1831 nand3_x0
xsubckt_731_oa22_x2 0 1542 1 291 357 553 oa22_x2
xsubckt_777_nor2_x0 1 0 1498 1499 1500 nor2_x0
xsubckt_848_nand2_x0 1 0 1437 1531 1799 nand2_x0
xsubckt_907_a2_x2 0 1388 1 1389 1391 a2_x2
xsubckt_1182_oa22_x2 0 1191 1 289 493 550 oa22_x2
xsubckt_1380_a4_x2 0 1020 1 1021 1033 1042 1051 a4_x2
xsubckt_1377_ao22_x2 0 1023 1 561 1138 1024 ao22_x2
xsubckt_563_o3_x2 0 116 1 287 466 587 o3_x2
xsubckt_351_nand2_x0 1 0 325 447 554 nand2_x0
xsubckt_300_nand3_x0 1 0 376 389 467 495 nand3_x0
xsubckt_654_nand4_x0 1 0 30 31 32 33 34 nand4_x0
xsubckt_997_a2_x2 0 1339 1 1340 1360 a2_x2
xsubckt_1883_sff1_x4 1 9 0 1601 1852 sff1_x4
xsubckt_1844_sff1_x4 1 9 0 1639 1765 sff1_x4
xsubckt_1805_sff1_x4 1 9 0 1670 1742 sff1_x4
xsubckt_1602_mx2_x2 0 804 1 978 805 838 mx2_x2
xsubckt_1601_mx2_x2 0 805 1 814 806 808 mx2_x2
xsubckt_1537_a3_x2 1 869 0 481 554 1771 a3_x2
xsubckt_1511_nand3_x0 1 0 895 904 920 961 nand3_x0
xsubckt_486_o2_x2 0 191 1 336 466 o2_x2
xsubckt_477_ao22_x2 0 200 1 533 515 527 ao22_x2
xsubckt_831_nand2_x0 1 0 1451 1520 1852 nand2_x0
xsubckt_968_nand2_x0 1 0 1680 1362 1363 nand2_x0
xsubckt_1068_a3_x2 1 1283 0 527 532 539 a3_x2
xsubckt_1082_nand2_x0 1 0 1270 1329 439 nand2_x0
xsubckt_1211_ao22_x2 0 1162 1 1180 1170 1163 ao22_x2
xsubckt_1263_a3_x2 1 1126 0 545 550 1865 a3_x2
xsubckt_1879_sff1_x4 1 9 0 1605 1775 sff1_x4
xsubckt_1642_ao22_x2 0 764 1 954 1540 1852 ao22_x2
xsubckt_1605_a2_x2 0 801 1 803 911 a2_x2
xsubckt_350_ao22_x2 0 326 1 434 327 328 ao22_x2
xsubckt_294_nand4_x0 1 0 382 1728 589 590 1729 nand4_x0
xsubckt_674_oa22_x2 0 12 1 281 360 630 oa22_x2
xsubckt_1047_oa22_x2 0 1665 1 1310 1309 1298 oa22_x2
xsubckt_1207_ao22_x2 0 1166 1 1726 382 322 ao22_x2
xsubckt_1791_sff1_x4 1 9 0 1684 1752 sff1_x4
xsubckt_1752_sff1_x4 1 9 0 1716 1842 sff1_x4
xsubckt_1292_nand2_x0 1 0 1100 1101 343 nand2_x0
xsubckt_414_nor4_x0 1 0 262 263 267 277 285 nor4_x0
xsubckt_647_nand3_x0 1 0 37 58 63 1828 nand3_x0
xsubckt_788_nand2_x0 1 0 1489 1543 1584 nand2_x0
xsubckt_1176_mx2_x2 0 1195 1 378 1196 1803 mx2_x2
xsubckt_1222_nor4_x0 1 0 1151 1152 1153 1156 1159 nor4_x0
xsubckt_1787_sff1_x4 1 9 0 1687 1783 sff1_x4
xsubckt_1685_a2_x2 0 721 1 723 730 a2_x2
xsubckt_1677_ao22_x2 0 729 1 735 737 940 ao22_x2
xsubckt_1347_nxr2_x1 1050 1 0 1053 1064 nxr2_x1
xsubckt_781_ao22_x2 0 1495 1 1527 1535 1850 ao22_x2
xsubckt_1024_nand2_x0 1 0 1314 438 623 nand2_x0
xsubckt_1061_nand3_x0 1 0 1288 1289 1336 1370 nand3_x0
xsubckt_1154_ao22_x2 0 1215 1 1216 1217 1218 ao22_x2
xsubckt_1177_mx2_x2 0 1638 1 1197 1195 1813 mx2_x2
xsubckt_1178_mx2_x2 0 1637 1 1721 1761 1883 mx2_x2
xsubckt_1704_nxr2_x1 702 1 0 703 795 nxr2_x1
xsubckt_1451_nand3_x0 1 0 954 325 360 377 nand3_x0
xsubckt_467_nand3_x0 1 0 210 481 495 556 nand3_x0
xsubckt_377_nand3_x0 1 0 299 404 409 525 nand3_x0
xsubckt_291_nand2_x0 1 0 385 387 1726 nand2_x0
xsubckt_720_nand3_x0 1 0 1552 57 63 1814 nand3_x0
xsubckt_771_nand2_x0 1 0 1905 1504 1510 nand2_x0
xsubckt_861_nand2_x0 1 0 1426 1520 1847 nand2_x0
xsubckt_1643_o2_x2 0 763 1 951 563 o2_x2
xsubckt_1546_ao22_x2 0 860 1 912 863 905 ao22_x2
xsubckt_1488_o2_x2 0 917 1 919 84 o2_x2
xsubckt_1361_nand3_x0 1 0 1038 545 550 1871 nand3_x0
xsubckt_630_nand3_x0 1 0 53 58 64 1845 nand3_x0
xsubckt_503_nand2_x0 1 0 175 177 255 nand2_x0
xsubckt_355_a4_x2 0 321 1 552 554 590 1729 a4_x2
xsubckt_335_a4_x2 0 341 1 342 344 348 350 a4_x2
xsubckt_1023_ao22_x2 0 1672 1 1325 1315 1319 ao22_x2
xsubckt_1493_ao22_x2 0 912 1 1523 461 1742 ao22_x2
xsubckt_590_a4_x2 0 91 1 286 290 374 376 a4_x2
xsubckt_450_nand3_x0 1 0 227 323 467 1726 nand3_x0
xsubckt_413_nand2_x0 1 0 263 264 265 nand2_x0
xsubckt_1144_nand2_x0 1 0 1642 1224 1226 nand2_x0
xsubckt_1271_nand3_x0 1 0 1119 358 554 666 nand3_x0
xsubckt_1583_nor3_x0 1 0 823 824 825 912 nor3_x0
xsubckt_1454_ao22_x2 0 951 1 553 480 309 ao22_x2
xsubckt_531_a2_x2 0 147 1 148 149 a2_x2
xsubckt_360_nand3_x0 1 0 316 447 1726 587 nand3_x0
xsubckt_336_a2_x2 0 340 1 341 352 a2_x2
xsubckt_737_a3_x2 1 1536 0 1537 1539 1541 a3_x2
xsubckt_840_nand3_x0 1 0 1444 1518 1526 1779 nand3_x0
xsubckt_891_nand2_x0 1 0 1401 1410 648 nand2_x0
xsubckt_932_a3_x2 1 1374 0 1414 57 64 a3_x2
xsubckt_981_nand2_x0 1 0 1676 1353 1354 nand2_x0
xsubckt_1216_oa22_x2 0 1157 1 494 492 480 oa22_x2
xsubckt_356_nand4_x0 1 0 320 552 554 590 1729 nand4_x0
xsubckt_158_ao22_x2 0 518 1 1786 1802 546 ao22_x2
xsubckt_105_inv_x0 1 0 564 1803 inv_x0
xsubckt_103_inv_x0 1 0 1790 565 inv_x0
xsubckt_102_inv_x0 1 0 1886 566 inv_x0
xsubckt_101_inv_x0 1 0 1807 567 inv_x0
xsubckt_100_inv_x0 1 0 1791 568 inv_x0
xsubckt_797_a3_x2 1 1481 0 1518 1526 1771 a3_x2
xsubckt_977_nand3_x0 1 0 1355 1365 406 412 nand3_x0
xsubckt_1003_a4_x2 0 1333 1 1336 1338 419 525 a4_x2
xsubckt_1608_oa22_x2 0 798 1 911 803 906 oa22_x2
xsubckt_109_inv_x0 1 0 562 1801 inv_x0
xsubckt_107_inv_x0 1 0 563 1802 inv_x0
xsubckt_246_o3_x2 0 430 1 431 468 471 o3_x2
xsubckt_712_oa22_x2 0 1559 1 48 482 643 oa22_x2
xsubckt_1073_a4_x2 0 1278 1 1292 173 525 539 a4_x2
xsubckt_480_nand3_x0 1 0 197 292 554 556 nand3_x0
xsubckt_139_o2_x2 0 537 1 1801 1786 o2_x2
xsubckt_302_nand3_x0 1 0 374 383 495 556 nand3_x0
xsubckt_910_mx2_x2 0 1385 1 355 1386 1798 mx2_x2
xsubckt_911_mx2_x2 0 1714 1 1413 1840 1385 mx2_x2
xsubckt_1083_a4_x2 0 1269 1 1272 1273 1329 439 a4_x2
xsubckt_1101_a3_x2 1 1255 0 1266 1292 520 a3_x2
xsubckt_1250_nand4_x0 1 0 1139 1140 1142 1534 185 nand4_x0
xsubckt_1864_sff1_x4 1 9 0 1620 1782 sff1_x4
xsubckt_1825_sff1_x4 1 9 0 1800 1808 sff1_x4
xsubckt_1715_ao22_x2 0 691 1 842 827 822 ao22_x2
xsubckt_1654_nand2_x0 1 0 752 754 756 nand2_x0
xsubckt_1620_a3_x2 1 786 0 481 554 1774 a3_x2
xsubckt_1513_nand3_x0 1 0 893 481 554 1770 nand3_x0
xsubckt_1424_nxr2_x1 980 1 0 981 989 nxr2_x1
xsubckt_1387_a4_x2 0 1014 1 1015 1016 1017 343 a4_x2
xsubckt_803_o2_x2 0 1475 1 1476 1481 o2_x2
xsubckt_833_nand2_x0 1 0 1891 1450 1454 nand2_x0
xsubckt_916_mx2_x2 0 1380 1 355 1381 1797 mx2_x2
xsubckt_917_mx2_x2 0 1713 1 1413 1839 1380 mx2_x2
xsubckt_1004_a2_x2 0 1332 1 1360 538 a2_x2
xsubckt_1171_a3_x2 1 1200 0 1201 1202 659 a3_x2
xsubckt_1500_o4_x2 0 905 1 911 918 919 84 o4_x2
xsubckt_1495_a3_x2 1 910 0 911 913 914 a3_x2
xsubckt_1416_mx2_x2 0 1606 1 656 988 1776 mx2_x2
xsubckt_1333_nand3_x0 1 0 1063 1065 1070 1078 nand3_x0
xsubckt_370_ao22_x2 0 306 1 662 441 307 ao22_x2
xsubckt_655_oa22_x2 0 1881 1 83 35 30 oa22_x2
xsubckt_780_nand3_x0 1 0 1496 1518 1526 1773 nand3_x0
xsubckt_1026_mx2_x2 0 1670 1 438 1318 1742 mx2_x2
xsubckt_1029_nand4_x0 1 0 1311 1312 173 401 413 nand4_x0
xsubckt_1772_sff1_x4 1 9 0 1702 1836 sff1_x4
xsubckt_1498_oa22_x2 0 907 1 961 920 910 oa22_x2
xsubckt_1378_a2_x2 0 1022 1 1023 1028 a2_x2
xsubckt_1371_mx2_x2 0 1610 1 656 1029 1780 mx2_x2
xsubckt_512_nand3_x0 1 0 166 404 410 525 nand3_x0
xsubckt_878_mx2_x2 0 1412 1 354 1803 1853 mx2_x2
xsubckt_879_mx2_x2 0 1719 1 1413 1845 1412 mx2_x2
xsubckt_1203_nor4_x0 1 0 1170 1171 1172 1190 1538 nor4_x0
xsubckt_1459_oa22_x2 0 946 1 1846 952 948 oa22_x2
xsubckt_596_nand4_x0 1 0 3 86 95 96 147 nand4_x0
xsubckt_21_inv_x0 1 0 1850 647 inv_x0
xsubckt_20_inv_x0 1 0 1851 648 inv_x0
xsubckt_920_nxr2_x1 1377 1 0 1378 1379 nxr2_x1
xsubckt_1768_sff1_x4 1 9 0 5 1727 sff1_x4
xsubckt_559_oa22_x2 0 120 1 170 174 436 oa22_x2
xsubckt_26_inv_x0 1 0 1846 642 inv_x0
xsubckt_25_inv_x0 1 0 1847 643 inv_x0
xsubckt_24_inv_x0 1 0 1855 644 inv_x0
xsubckt_23_inv_x0 1 0 1848 645 inv_x0
xsubckt_22_inv_x0 1 0 1849 646 inv_x0
xsubckt_863_nand2_x0 1 0 1900 1425 1429 nand2_x0
xsubckt_1566_ao22_x2 0 840 1 560 951 1016 ao22_x2
xsubckt_126_a3_x2 1 550 0 551 552 554 a3_x2
xsubckt_29_inv_x0 1 0 1765 639 inv_x0
xsubckt_28_inv_x0 1 0 1754 640 inv_x0
xsubckt_27_inv_x0 1 0 1757 641 inv_x0
xsubckt_238_nand4_x0 1 0 438 551 552 554 1721 nand4_x0
xsubckt_293_a4_x2 0 383 1 1728 589 590 1729 a4_x2
xsubckt_1043_ao22_x2 0 1300 1 507 511 1812 ao22_x2
xsubckt_587_a4_x2 0 94 1 220 221 272 276 a4_x2
xsubckt_577_a4_x2 0 103 1 330 333 455 458 a4_x2
xsubckt_567_a4_x2 0 112 1 113 120 121 142 a4_x2
xsubckt_1536_nand2_x0 1 0 870 872 885 nand2_x0
xsubckt_325_nand2_x0 1 0 351 362 495 nand2_x0
xsubckt_214_a2_x2 0 462 1 463 465 a2_x2
xsubckt_805_nand2_x0 1 0 1474 1543 1561 nand2_x0
xsubckt_850_a3_x2 1 1435 0 1436 1437 1438 a3_x2
xsubckt_898_nxr2_x1 1395 1 0 1396 1397 nxr2_x1
xsubckt_1446_nand2_x0 1 0 959 1189 334 nand2_x0
xsubckt_274_a2_x2 0 402 1 526 532 a2_x2
xsubckt_743_nor2_x0 1 0 1530 269 449 nor2_x0
xsubckt_880_a3_x2 1 1411 0 1854 1764 1762 a3_x2
xsubckt_1410_a4_x2 0 993 1 994 995 996 343 a4_x2
xsubckt_1356_nand2_x0 1 0 1042 1044 1049 nand2_x0
xsubckt_1304_ao22_x2 0 1089 1 629 1129 1091 ao22_x2
xsubckt_588_a2_x2 0 93 1 94 114 a2_x2
xsubckt_418_o3_x2 0 8 1 259 391 396 o3_x2
xsubckt_793_a2_x2 0 1484 1 1485 1486 a2_x2
xsubckt_1089_nand4_x0 1 0 1264 1326 173 525 539 nand4_x0
xsubckt_1810_sff1_x4 1 9 0 1665 1734 sff1_x4
xsubckt_728_oa22_x2 0 1875 1 83 1550 1545 oa22_x2
xsubckt_767_oa22_x2 0 1507 1 1521 1522 610 oa22_x2
xsubckt_1125_nand3_x0 1 0 1241 1419 654 658 nand3_x0
xsubckt_1884_sff1_x4 1 9 0 1600 1851 sff1_x4
xsubckt_1693_nand3_x0 1 0 713 714 717 720 nand3_x0
xsubckt_1612_mx2_x2 0 794 1 804 798 800 mx2_x2
xsubckt_1611_mx2_x2 0 795 1 804 799 801 mx2_x2
xsubckt_1515_nand3_x0 1 0 891 932 937 1797 nand3_x0
xsubckt_1290_ao22_x2 0 1102 1 1130 372 1773 ao22_x2
xsubckt_533_nor3_x0 1 0 145 1724 1855 1723 nor3_x0
xsubckt_392_nand3_x0 1 0 284 292 467 493 nand3_x0
xsubckt_711_o2_x2 0 1560 1 51 613 o2_x2
xsubckt_835_nand2_x0 1 0 1448 1458 1871 nand2_x0
xsubckt_1035_nand3_x0 1 0 1307 407 505 515 nand3_x0
xsubckt_1086_nand2_x0 1 0 1267 438 583 nand2_x0
xsubckt_1098_nor2_x0 1 0 1655 1257 1261 nor2_x0
xsubckt_1212_ao22_x2 0 1161 1 362 481 495 ao22_x2
xsubckt_1845_sff1_x4 1 9 0 1638 1813 sff1_x4
xsubckt_1806_sff1_x4 1 9 0 1669 1738 sff1_x4
xsubckt_636_oa22_x2 0 47 1 337 484 494 oa22_x2
xsubckt_439_ao22_x2 0 238 1 338 473 495 ao22_x2
xsubckt_1206_a2_x2 0 1167 1 1169 1534 a2_x2
xsubckt_1247_ao22_x2 0 1142 1 549 545 496 ao22_x2
xsubckt_1256_a2_x2 0 1133 1 1134 549 a2_x2
xsubckt_1792_sff1_x4 1 9 0 1683 1740 sff1_x4
xsubckt_1753_sff1_x4 1 9 0 1715 1841 sff1_x4
xsubckt_1735_a2_x2 0 672 1 673 713 a2_x2
xsubckt_1391_nxr2_x1 1010 1 0 1012 1020 nxr2_x1
xsubckt_1386_nand2_x0 1 0 1015 372 1849 nand2_x0
xsubckt_551_nand4_x0 1 0 128 275 467 586 1725 nand4_x0
xsubckt_1229_mx2_x2 0 1636 1 1145 1906 1865 mx2_x2
xsubckt_1576_mx2_x2 0 830 1 833 927 940 mx2_x2
xsubckt_598_nand4_x0 1 0 84 85 281 356 360 nand4_x0
xsubckt_334_nand3_x0 1 0 342 358 554 556 nand3_x0
xsubckt_904_nand3_x0 1 0 1391 1855 1764 1762 nand3_x0
xsubckt_955_nand2_x0 1 0 1371 438 1740 nand2_x0
xsubckt_1014_nand4_x0 1 0 1322 419 504 517 520 nand4_x0
xsubckt_1788_sff1_x4 1 9 0 1722 1784 sff1_x4
xsubckt_1749_sff1_x4 1 9 0 1719 1845 sff1_x4
xsubckt_1686_nand2_x0 1 0 720 723 730 nand2_x0
xsubckt_1639_ao22_x2 0 767 1 912 770 905 ao22_x2
xsubckt_1590_ao22_x2 0 816 1 647 953 818 ao22_x2
xsubckt_1551_ao22_x2 0 855 1 645 953 857 ao22_x2
xsubckt_1313_oa22_x2 0 1081 1 1848 1135 1083 oa22_x2
xsubckt_295_nand2_x0 1 0 381 383 493 nand2_x0
xsubckt_775_nand2_x0 1 0 1500 1501 1502 nand2_x0
xsubckt_865_nand2_x0 1 0 1423 1458 1866 nand2_x0
xsubckt_1065_nand3_x0 1 0 1285 1286 203 512 nand3_x0
xsubckt_1705_nxr2_x1 701 1 0 703 794 nxr2_x1
xsubckt_1548_o2_x2 0 858 1 951 559 o2_x2
xsubckt_1508_o2_x2 0 898 1 899 901 o2_x2
xsubckt_544_nand3_x0 1 0 6 135 151 162 nand3_x0
xsubckt_513_a3_x2 1 165 0 166 167 168 a3_x2
xsubckt_338_a3_x2 1 338 0 490 590 1729 a3_x2
xsubckt_660_a4_x2 0 25 1 26 27 28 29 a4_x2
xsubckt_709_a4_x2 0 1562 1 1563 1564 1565 1566 a4_x2
xsubckt_1267_nor2_x0 1 0 1122 1123 1124 nor2_x0
xsubckt_608_ao22_x2 0 75 1 586 322 287 ao22_x2
xsubckt_583_a3_x2 1 97 0 98 99 129 a3_x2
xsubckt_543_a3_x2 1 135 0 136 392 397 a3_x2
xsubckt_132_a2_x2 0 544 1 565 1786 a2_x2
xsubckt_223_nand4_x0 1 0 453 490 587 1730 591 nand4_x0
xsubckt_807_nand2_x0 1 0 1472 1525 1847 nand2_x0
xsubckt_1007_nand3_x0 1 0 1329 1331 173 525 nand3_x0
xsubckt_1311_nand2_x0 1 0 1083 1085 343 nand2_x0
xsubckt_613_nand4_x0 1 0 70 71 77 549 1731 nand4_x0
xsubckt_476_a2_x2 0 201 1 202 204 a2_x2
xsubckt_400_nand2_x0 1 0 276 449 467 nand2_x0
xsubckt_111_inv_x0 1 0 561 1800 inv_x0
xsubckt_703_nand4_x0 1 0 1567 1568 1569 1570 43 nand4_x0
xsubckt_877_a3_x2 1 1413 0 1414 58 64 a3_x2
xsubckt_1095_nand3_x0 1 0 1259 1294 1338 525 nand3_x0
xsubckt_1648_oa22_x2 0 758 1 35 956 760 oa22_x2
xsubckt_1560_oa22_x2 0 846 1 849 850 926 oa22_x2
xsubckt_1395_nand3_x0 1 0 1007 545 550 1868 nand3_x0
xsubckt_1324_ao22_x2 0 1071 1 627 1129 1073 ao22_x2
xsubckt_574_nand3_x0 1 0 105 106 109 427 nand3_x0
xsubckt_496_a2_x2 0 182 1 183 299 a2_x2
xsubckt_117_inv_x0 1 0 558 1797 inv_x0
xsubckt_115_inv_x0 1 0 559 1798 inv_x0
xsubckt_113_inv_x0 1 0 560 1799 inv_x0
xsubckt_249_nor3_x0 1 0 427 428 433 440 nor3_x0
xsubckt_713_oa22_x2 0 1558 1 281 360 627 oa22_x2
xsubckt_791_oa22_x2 0 1486 1 1521 1522 607 oa22_x2
xsubckt_1131_nand2_x0 1 0 1235 549 1797 nand2_x0
xsubckt_1830_sff1_x4 1 9 0 1653 1746 sff1_x4
xsubckt_1521_nand2_x0 1 0 885 887 905 nand2_x0
xsubckt_484_nand3_x0 1 0 193 489 495 556 nand3_x0
xsubckt_447_nand2_x0 1 0 230 232 405 nand2_x0
xsubckt_119_inv_x0 1 0 557 1796 inv_x0
xsubckt_787_oa22_x2 0 1897 1 13 1543 1490 oa22_x2
xsubckt_921_mx2_x2 0 1376 1 355 1377 1796 mx2_x2
xsubckt_1254_nand4_x0 1 0 1135 1534 369 385 491 nand4_x0
xsubckt_1556_oa22_x2 0 850 1 866 868 939 oa22_x2
xsubckt_1517_oa22_x2 0 889 1 891 893 916 oa22_x2
xsubckt_1341_nand2_x0 1 0 1056 372 1853 nand2_x0
xsubckt_610_nand2_x0 1 0 73 316 345 nand2_x0
xsubckt_424_ao22_x2 0 253 1 436 254 258 ao22_x2
xsubckt_259_o2_x2 0 417 1 1798 1786 o2_x2
xsubckt_837_nand2_x0 1 0 1446 1531 1801 nand2_x0
xsubckt_922_mx2_x2 0 1712 1 1413 1838 1376 mx2_x2
xsubckt_924_mx2_x2 0 1711 1 1375 1821 1412 mx2_x2
xsubckt_925_mx2_x2 0 1710 1 1375 1820 1403 mx2_x2
xsubckt_926_mx2_x2 0 1709 1 1375 1819 1398 mx2_x2
xsubckt_927_mx2_x2 0 1708 1 1375 1818 1394 mx2_x2
xsubckt_964_nand3_x0 1 0 1364 1365 150 412 nand3_x0
xsubckt_1072_oa22_x2 0 1279 1 1280 1282 403 oa22_x2
xsubckt_1074_nand4_x0 1 0 1277 1292 173 525 539 nand4_x0
xsubckt_1251_a3_x2 1 1138 0 1534 385 491 a3_x2
xsubckt_1865_sff1_x4 1 9 0 1619 1781 sff1_x4
xsubckt_1826_sff1_x4 1 9 0 1799 1807 sff1_x4
xsubckt_1425_mx2_x2 0 1605 1 656 980 1775 mx2_x2
xsubckt_748_o2_x2 0 1525 1 1527 1535 o2_x2
xsubckt_928_mx2_x2 0 1707 1 1375 1817 1393 mx2_x2
xsubckt_929_mx2_x2 0 1706 1 1375 1816 1385 mx2_x2
xsubckt_1033_mx2_x2 0 1668 1 438 1345 1733 mx2_x2
xsubckt_1164_a2_x2 0 1206 1 1207 1208 a2_x2
xsubckt_1174_a2_x2 0 1197 1 1198 1199 a2_x2
xsubckt_1653_a2_x2 0 753 1 754 756 a2_x2
xsubckt_1641_nand2_x0 1 0 765 766 773 nand2_x0
xsubckt_1382_mx2_x2 0 1609 1 656 1019 1779 mx2_x2
xsubckt_694_nand3_x0 1 0 1576 57 64 1832 nand3_x0
xsubckt_888_mx2_x2 0 1403 1 355 1404 1802 mx2_x2
xsubckt_889_mx2_x2 0 1718 1 1413 1844 1403 mx2_x2
xsubckt_1161_nand2_x0 1 0 1209 1210 482 nand2_x0
xsubckt_1194_a2_x2 0 1179 1 79 369 a2_x2
xsubckt_1773_sff1_x4 1 9 0 1701 1835 sff1_x4
xsubckt_1673_a2_x2 0 733 1 734 736 a2_x2
xsubckt_1478_a2_x2 0 927 1 928 941 a2_x2
xsubckt_906_nand3_x0 1 0 1389 644 650 1762 nand3_x0
xsubckt_1102_o2_x2 0 1254 1 1255 1278 o2_x2
xsubckt_1769_sff1_x4 1 9 0 4 1726 sff1_x4
xsubckt_160_nand2_x0 1 0 516 518 519 nand2_x0
xsubckt_33_inv_x0 1 0 1747 635 inv_x0
xsubckt_32_inv_x0 1 0 1785 636 inv_x0
xsubckt_31_inv_x0 1 0 1766 637 inv_x0
xsubckt_30_inv_x0 1 0 1813 638 inv_x0
xsubckt_297_nand2_x0 1 0 379 380 384 nand2_x0
xsubckt_867_nand2_x0 1 0 1421 1520 1846 nand2_x0
xsubckt_353_a4_x2 0 323 1 552 587 590 1729 a4_x2
xsubckt_39_inv_x0 1 0 1772 629 inv_x0
xsubckt_38_inv_x0 1 0 1773 630 inv_x0
xsubckt_37_inv_x0 1 0 1774 631 inv_x0
xsubckt_36_inv_x0 1 0 1781 632 inv_x0
xsubckt_35_inv_x0 1 0 1782 633 inv_x0
xsubckt_34_inv_x0 1 0 1738 634 inv_x0
xsubckt_673_nand4_x0 1 0 13 15 16 17 18 nand4_x0
xsubckt_798_ao22_x2 0 1480 1 1527 1535 1848 ao22_x2
xsubckt_1103_nand2_x0 1 0 1253 1335 515 nand2_x0
xsubckt_1725_oa22_x2 0 681 1 682 895 908 oa22_x2
xsubckt_1567_ao22_x2 0 839 1 646 953 840 ao22_x2
xsubckt_1528_ao22_x2 0 878 1 892 894 940 ao22_x2
xsubckt_632_ao22_x2 0 51 1 492 357 279 ao22_x2
xsubckt_456_nand3_x0 1 0 221 467 485 495 nand3_x0
xsubckt_433_oa22_x2 0 244 1 493 292 346 oa22_x2
xsubckt_198_a4_x2 0 478 1 479 482 486 491 a4_x2
xsubckt_1191_nand2_x0 1 0 1182 1186 1188 nand2_x0
xsubckt_1276_nxr2_x1 1114 1 0 1116 1124 nxr2_x1
xsubckt_1530_nand3_x0 1 0 876 891 893 927 nand3_x0
xsubckt_471_a3_x2 1 206 0 207 217 224 a3_x2
xsubckt_461_a3_x2 1 216 0 481 554 556 a3_x2
xsubckt_324_a2_x2 0 352 1 353 359 a2_x2
xsubckt_190_nand2_x0 1 0 486 489 493 nand2_x0
xsubckt_760_nand2_x0 1 0 1513 1514 1515 nand2_x0
xsubckt_846_nand3_x0 1 0 1439 1518 1526 1778 nand3_x0
xsubckt_1009_nand3_x0 1 0 1327 1328 1329 439 nand3_x0
xsubckt_1169_nor3_x0 1 0 1202 1755 1763 1734 nor3_x0
xsubckt_1350_nand3_x0 1 0 1048 545 550 1872 nand3_x0
xsubckt_364_a2_x2 0 312 1 313 315 a2_x2
xsubckt_344_a2_x2 0 332 1 338 493 a2_x2
xsubckt_159_a2_x2 0 517 1 518 519 a2_x2
xsubckt_149_a2_x2 0 527 1 529 531 a2_x2
xsubckt_756_nand3_x0 1 0 1517 1518 1526 1782 nand3_x0
xsubckt_970_a3_x2 1 1360 0 420 506 509 a3_x2
xsubckt_1309_nand3_x0 1 0 1085 545 550 1860 nand3_x0
xsubckt_873_a2_x2 0 1417 1 1419 1746 a2_x2
xsubckt_1051_a4_x2 0 1295 1 439 517 520 533 a4_x2
xsubckt_1650_nand3_x0 1 0 756 481 554 1781 nand3_x0
xsubckt_1850_sff1_x4 1 9 0 1634 1863 sff1_x4
xsubckt_1811_sff1_x4 1 9 0 1664 1763 sff1_x4
xsubckt_1519_nand3_x0 1 0 887 889 890 911 nand3_x0
xsubckt_1433_nand2_x0 1 0 972 461 1755 nand2_x0
xsubckt_396_nand3_x0 1 0 280 292 467 554 nand3_x0
xsubckt_218_nand3_x0 1 0 458 467 493 499 nand3_x0
xsubckt_641_oa22_x2 0 42 1 44 343 638 oa22_x2
xsubckt_768_oa22_x2 0 1506 1 331 446 563 oa22_x2
xsubckt_790_nand2_x0 1 0 1487 1525 1849 nand2_x0
xsubckt_839_nand2_x0 1 0 1904 1445 1449 nand2_x0
xsubckt_1248_a3_x2 1 1141 0 266 345 386 a3_x2
xsubckt_1885_sff1_x4 1 9 0 1599 1850 sff1_x4
xsubckt_1846_sff1_x4 1 9 0 1592 1762 sff1_x4
xsubckt_1807_sff1_x4 1 9 0 1668 1733 sff1_x4
xsubckt_1473_a3_x2 1 932 0 933 934 936 a3_x2
xsubckt_125_nor2_x0 1 0 551 1730 1729 nor2_x0
xsubckt_686_o2_x2 0 1583 1 51 615 o2_x2
xsubckt_1052_a2_x2 0 1294 1 1360 413 a2_x2
xsubckt_1230_mx2_x2 0 1635 1 1145 1905 1864 mx2_x2
xsubckt_1231_mx2_x2 0 1634 1 1145 1898 1863 mx2_x2
xsubckt_1232_mx2_x2 0 1633 1 1145 1897 1862 mx2_x2
xsubckt_1233_mx2_x2 0 1632 1 1145 1896 1861 mx2_x2
xsubckt_1628_mx2_x2 0 778 1 781 927 940 mx2_x2
xsubckt_1541_a2_x2 0 865 1 866 868 a2_x2
xsubckt_1445_oa22_x2 0 960 1 495 489 323 oa22_x2
xsubckt_1339_nand3_x0 1 0 1058 545 550 1873 nand3_x0
xsubckt_569_nor3_x0 1 0 110 194 277 285 nor3_x0
xsubckt_518_nand3_x0 1 0 160 362 495 556 nand3_x0
xsubckt_676_oa22_x2 0 10 1 48 482 647 oa22_x2
xsubckt_696_nand3_x0 1 0 1574 57 63 1816 nand3_x0
xsubckt_1092_a2_x2 0 1656 1 1262 1267 a2_x2
xsubckt_1158_o4_x2 0 1212 1 1217 1418 1760 1755 o4_x2
xsubckt_1234_mx2_x2 0 1631 1 1145 1895 1860 mx2_x2
xsubckt_1235_mx2_x2 0 1630 1 1145 1894 1859 mx2_x2
xsubckt_1236_mx2_x2 0 1629 1 1145 1893 1858 mx2_x2
xsubckt_1237_mx2_x2 0 1628 1 1145 1892 1873 mx2_x2
xsubckt_1238_mx2_x2 0 1627 1 1145 1891 1872 mx2_x2
xsubckt_1239_mx2_x2 0 1626 1 1145 1904 1871 mx2_x2
xsubckt_1793_sff1_x4 1 9 0 1682 1741 sff1_x4
xsubckt_1754_sff1_x4 1 9 0 1714 1840 sff1_x4
xsubckt_506_nxr2_x1 172 1 0 517 520 nxr2_x1
xsubckt_201_nand3_x0 1 0 475 476 490 586 nand3_x0
xsubckt_822_nand2_x0 1 0 1459 1531 1803 nand2_x0
xsubckt_1789_sff1_x4 1 9 0 1686 1754 sff1_x4
xsubckt_1710_nxr2_x1 696 1 0 704 707 nxr2_x1
xsubckt_162_nand2_x0 1 0 514 516 521 nand2_x0
xsubckt_299_nand2_x0 1 0 377 389 495 nand2_x0
xsubckt_869_nand2_x0 1 0 1899 1420 1424 nand2_x0
xsubckt_552_nand2_x0 1 0 127 317 556 nand2_x0
xsubckt_271_a4_x2 0 405 1 412 420 504 538 a4_x2
xsubckt_1460_ao22_x2 0 945 1 1551 957 947 ao22_x2
xsubckt_1025_ao22_x2 0 1671 1 1325 1320 1314 ao22_x2
xsubckt_1193_nor3_x0 1 0 1180 1182 1183 1190 nor3_x0
xsubckt_1279_nand3_x0 1 0 1112 545 550 1863 nand3_x0
xsubckt_623_a3_x2 1 60 0 61 71 77 a3_x2
xsubckt_595_a4_x2 0 86 1 87 90 133 326 a4_x2
xsubckt_428_a3_x2 1 249 0 251 504 538 a3_x2
xsubckt_762_nand2_x0 1 0 1511 1512 1517 nand2_x0
xsubckt_1456_ao22_x2 0 949 1 557 951 984 ao22_x2
xsubckt_1352_nand3_x0 1 0 1046 383 554 1872 nand3_x0
xsubckt_272_a2_x2 0 404 1 516 520 a2_x2
xsubckt_576_a2_x2 0 104 1 117 253 a2_x2
xsubckt_556_a2_x2 0 123 1 124 126 a2_x2
xsubckt_492_nand2_x0 1 0 7 186 205 nand2_x0
xsubckt_188_nand3_x0 1 0 488 490 1730 591 nand3_x0
xsubckt_668_nand3_x0 1 0 18 57 63 1818 nand3_x0
xsubckt_751_a2_x2 0 1522 1 1524 482 a2_x2
xsubckt_792_oa22_x2 0 1485 1 331 446 560 oa22_x2
xsubckt_987_a3_x2 1 1348 0 256 404 533 a3_x2
xsubckt_1652_nand3_x0 1 0 754 932 937 1802 nand3_x0
xsubckt_1615_nand2_x0 1 0 791 792 1037 nand2_x0
xsubckt_1525_nand2_x0 1 0 881 883 884 nand2_x0
xsubckt_1522_oa22_x2 0 884 1 955 1541 643 oa22_x2
xsubckt_210_o2_x2 0 466 1 2 1721 o2_x2
xsubckt_714_oa22_x2 0 1557 1 44 343 637 oa22_x2
xsubckt_972_nand2_x0 1 0 1679 1359 1361 nand2_x0
xsubckt_1038_a4_x2 0 1305 1 551 554 1727 1721 a4_x2
xsubckt_1045_nand2_x0 1 0 1666 1299 1303 nand2_x0
xsubckt_1172_nand3_x0 1 0 1199 485 495 1734 nand3_x0
xsubckt_1253_a4_x2 0 1136 1 1534 369 385 491 a4_x2
xsubckt_1870_sff1_x4 1 9 0 1614 1770 sff1_x4
xsubckt_1831_sff1_x4 1 9 0 1652 1786 sff1_x4
xsubckt_1721_ao22_x2 0 685 1 687 688 843 ao22_x2
xsubckt_1489_nor3_x0 1 0 916 918 919 84 nor3_x0
xsubckt_1435_nand2_x0 1 0 970 971 1523 nand2_x0
xsubckt_930_mx2_x2 0 1705 1 1375 1815 1380 mx2_x2
xsubckt_931_mx2_x2 0 1704 1 1375 1814 1376 mx2_x2
xsubckt_933_mx2_x2 0 1703 1 1374 1837 1412 mx2_x2
xsubckt_934_mx2_x2 0 1702 1 1374 1836 1403 mx2_x2
xsubckt_1168_nand4_x0 1 0 1203 551 552 554 662 nand4_x0
xsubckt_1866_sff1_x4 1 9 0 1618 1774 sff1_x4
xsubckt_1562_mx3_x2 1 0 844 977 852 880 847 850 mx3_x2
xsubckt_1561_mx3_x2 1 0 845 977 852 879 846 851 mx3_x2
xsubckt_1345_nand2_x0 1 0 1052 1054 1060 nand2_x0
xsubckt_561_nand3_x0 1 0 118 232 249 437 nand3_x0
xsubckt_401_nor4_x0 1 0 275 1728 1727 1730 1729 nor4_x0
xsubckt_935_mx2_x2 0 1701 1 1374 1835 1398 mx2_x2
xsubckt_936_mx2_x2 0 1700 1 1374 1834 1394 mx2_x2
xsubckt_937_mx2_x2 0 1699 1 1374 1833 1393 mx2_x2
xsubckt_938_mx2_x2 0 1698 1 1374 1832 1385 mx2_x2
xsubckt_939_mx2_x2 0 1697 1 1374 1831 1380 mx2_x2
xsubckt_1196_a3_x2 1 1177 0 375 381 482 a3_x2
xsubckt_1827_sff1_x4 1 9 0 1798 1806 sff1_x4
xsubckt_434_nand2_x0 1 0 243 432 478 nand2_x0
xsubckt_894_mx2_x2 0 1398 1 355 1399 1801 mx2_x2
xsubckt_895_mx2_x2 0 1717 1 1413 1843 1398 mx2_x2
xsubckt_1114_nand3_x0 1 0 1652 1244 193 313 nand3_x0
xsubckt_1151_nand4_x0 1 0 1218 1243 377 482 549 nand4_x0
xsubckt_1175_mx3_x2 1 0 1196 1202 1740 1855 1853 661 mx3_x2
xsubckt_1274_a2_x2 0 1116 1 1117 1121 a2_x2
xsubckt_1774_sff1_x4 1 9 0 1700 1834 sff1_x4
xsubckt_1392_mx2_x2 0 1608 1 656 1010 1778 mx2_x2
xsubckt_381_nand3_x0 1 0 295 402 404 539 nand3_x0
xsubckt_824_nand2_x0 1 0 1457 1458 1873 nand2_x0
xsubckt_899_mx2_x2 0 1394 1 355 1395 1800 mx2_x2
xsubckt_1048_mx2_x2 0 1664 1 1304 1302 1763 mx2_x2
xsubckt_1730_nxr2_x1 676 1 0 683 685 nxr2_x1
xsubckt_1699_ao22_x2 0 707 1 710 712 738 ao22_x2
xsubckt_1334_oa22_x2 0 1062 1 1078 1070 1065 oa22_x2
xsubckt_40_inv_x0 1 0 1771 628 inv_x0
xsubckt_241_ao22_x2 0 435 1 544 540 437 ao22_x2
xsubckt_681_nand3_x0 1 0 1588 57 63 1817 nand3_x0
xsubckt_1726_nxr2_x1 680 1 0 681 896 nxr2_x1
xsubckt_1506_o2_x2 0 900 1 951 564 o2_x2
xsubckt_41_inv_x0 1 0 1770 627 inv_x0
xsubckt_42_inv_x0 1 0 1769 626 inv_x0
xsubckt_43_inv_x0 1 0 1745 625 inv_x0
xsubckt_44_inv_x0 1 0 1744 624 inv_x0
xsubckt_45_inv_x0 1 0 1743 623 inv_x0
xsubckt_46_inv_x0 1 0 1742 622 inv_x0
xsubckt_1266_nor3_x0 1 0 1123 1125 1127 1139 nor3_x0
xsubckt_1675_nand2_x0 1 0 731 732 911 nand2_x0
xsubckt_1568_ao22_x2 0 838 1 1585 957 839 ao22_x2
xsubckt_1369_oa22_x2 0 1030 1 1051 1042 1033 oa22_x2
xsubckt_409_nand4_x0 1 0 267 268 271 272 276 nand4_x0
xsubckt_374_nand2_x0 1 0 302 489 495 nand2_x0
xsubckt_323_nand3_x0 1 0 353 358 493 556 nand3_x0
xsubckt_47_inv_x0 1 0 1741 621 inv_x0
xsubckt_48_inv_x0 1 0 1768 620 inv_x0
xsubckt_49_inv_x0 1 0 1767 619 inv_x0
xsubckt_1054_nand3_x0 1 0 1663 1293 1296 1297 nand3_x0
xsubckt_1645_nor2_x0 1 0 761 762 764 nor2_x0
xsubckt_1585_nand2_x0 1 0 821 822 905 nand2_x0
xsubckt_571_a3_x2 1 108 0 113 217 224 a3_x2
xsubckt_541_a3_x2 1 137 0 138 293 363 a3_x2
xsubckt_521_a3_x2 1 157 0 158 159 160 a3_x2
xsubckt_376_a3_x2 1 300 0 404 409 525 a3_x2
xsubckt_120_a2_x2 0 556 1 655 1721 a2_x2
xsubckt_233_nand3_x0 1 0 443 445 446 452 nand3_x0
xsubckt_319_nand4_x0 1 0 357 588 1727 590 1729 nand4_x0
xsubckt_764_nand2_x0 1 0 1510 1543 35 nand2_x0
xsubckt_854_nand2_x0 1 0 1432 1520 1848 nand2_x0
xsubckt_591_a3_x2 1 90 0 91 92 93 a3_x2
xsubckt_581_a3_x2 1 99 0 100 101 139 a3_x2
xsubckt_180_nand4_x0 1 0 496 552 586 1730 591 nand4_x0
xsubckt_194_nand2_x0 1 0 482 485 495 nand2_x0
xsubckt_239_a2_x2 0 437 1 439 655 a2_x2
xsubckt_1707_nand2_x0 1 0 699 461 1764 nand2_x0
xsubckt_1542_nxr2_x1 864 1 0 865 915 nxr2_x1
xsubckt_443_nand3_x0 1 0 234 383 467 493 nand3_x0
xsubckt_406_nand2_x0 1 0 270 275 587 nand2_x0
xsubckt_279_a2_x2 0 397 1 398 423 a2_x2
xsubckt_316_nand2_x0 1 0 360 362 493 nand2_x0
xsubckt_913_a2_x2 0 1383 1 1391 643 a2_x2
xsubckt_1503_oa22_x2 0 1604 1 903 907 979 oa22_x2
xsubckt_1448_nor4_x0 1 0 957 958 959 1172 76 nor4_x0
xsubckt_207_o2_x2 0 469 1 1724 1855 o2_x2
xsubckt_212_nand4_x0 1 0 464 551 552 586 1725 nand4_x0
xsubckt_226_nand2_x0 1 0 450 1726 1725 nand2_x0
xsubckt_773_oa22_x2 0 1502 1 1521 1522 609 oa22_x2
xsubckt_1084_nand3_x0 1 0 1268 1269 1279 1334 nand3_x0
xsubckt_1181_a4_x2 0 1192 1 551 587 1728 589 a4_x2
xsubckt_1890_sff1_x4 1 9 0 1594 1854 sff1_x4
xsubckt_1851_sff1_x4 1 9 0 1633 1862 sff1_x4
xsubckt_1812_sff1_x4 1 9 0 1663 1749 sff1_x4
xsubckt_1474_nand3_x0 1 0 931 932 937 1796 nand3_x0
xsubckt_412_o2_x2 0 264 1 452 466 o2_x2
xsubckt_1886_sff1_x4 1 9 0 1598 1849 sff1_x4
xsubckt_1632_mx2_x2 0 774 1 788 776 780 mx2_x2
xsubckt_1631_mx2_x2 0 775 1 788 777 779 mx2_x2
xsubckt_1384_nand3_x0 1 0 1017 545 550 1869 nand3_x0
xsubckt_165_nor2_x0 1 0 511 1796 1786 nor2_x0
xsubckt_690_nand4_x0 1 0 1579 1580 1581 1583 44 nand4_x0
xsubckt_726_o2_x2 0 1546 1 51 612 o2_x2
xsubckt_1112_a2_x2 0 1245 1 655 1786 a2_x2
xsubckt_1132_a2_x2 0 1234 1 1847 1740 a2_x2
xsubckt_1240_mx2_x2 0 1625 1 1145 1903 1870 mx2_x2
xsubckt_1257_nand2_x0 1 0 1132 1134 549 nand2_x0
xsubckt_1847_sff1_x4 1 9 0 1637 1761 sff1_x4
xsubckt_1808_sff1_x4 1 9 0 1667 1755 sff1_x4
xsubckt_1634_mx2_x2 0 772 1 978 775 814 mx2_x2
xsubckt_1633_mx2_x2 0 773 1 978 774 813 mx2_x2
xsubckt_1426_a2_x2 0 979 1 1856 656 a2_x2
xsubckt_638_oa22_x2 0 45 1 48 482 652 oa22_x2
xsubckt_473_nand3_x0 1 0 204 338 467 493 nand3_x0
xsubckt_436_nand2_x0 1 0 241 338 495 nand2_x0
xsubckt_422_nand4_x0 1 0 255 413 419 504 538 nand4_x0
xsubckt_649_nand4_x0 1 0 35 37 38 39 40 nand4_x0
xsubckt_677_oa22_x2 0 1591 1 44 343 665 oa22_x2
xsubckt_1241_mx2_x2 0 1624 1 1145 1902 1869 mx2_x2
xsubckt_1242_mx2_x2 0 1623 1 1145 1901 1868 mx2_x2
xsubckt_1243_mx2_x2 0 1622 1 1145 1900 1867 mx2_x2
xsubckt_1244_mx2_x2 0 1621 1 1145 1899 1866 mx2_x2
xsubckt_1794_sff1_x4 1 9 0 1681 1759 sff1_x4
xsubckt_1755_sff1_x4 1 9 0 1713 1839 sff1_x4
xsubckt_1691_a2_x2 0 715 1 722 731 a2_x2
xsubckt_1681_a2_x2 0 725 1 726 925 a2_x2
xsubckt_722_nand4_x0 1 0 1550 1552 1553 1554 1555 nand4_x0
xsubckt_1711_nxr2_x1 695 1 0 704 706 nxr2_x1
xsubckt_1599_mx2_x2 0 807 1 809 927 940 mx2_x2
xsubckt_1594_nand3_x0 1 0 812 481 554 1773 nand3_x0
xsubckt_683_nand3_x0 1 0 1586 57 64 1833 nand3_x0
xsubckt_1630_nand2_x0 1 0 776 778 925 nand2_x0
xsubckt_1592_ao22_x2 0 814 1 14 957 816 ao22_x2
xsubckt_1553_ao22_x2 0 853 1 1572 957 855 ao22_x2
xsubckt_1315_oa22_x2 0 1079 1 1771 1128 1081 oa22_x2
xsubckt_199_nand4_x0 1 0 477 479 482 486 491 nand4_x0
xsubckt_1588_ao22_x2 0 818 1 561 951 1025 ao22_x2
xsubckt_1549_ao22_x2 0 857 1 559 951 1006 ao22_x2
xsubckt_1297_nxr2_x1 1095 1 0 1098 1106 nxr2_x1
xsubckt_452_nand4_x0 1 0 225 257 404 437 525 nand4_x0
xsubckt_1422_ao22_x2 0 982 1 557 1138 983 ao22_x2
xsubckt_1360_nand2_x0 1 0 1039 1137 1801 nand2_x0
xsubckt_130_ao22_x2 0 546 1 1795 616 664 ao22_x2
xsubckt_244_a3_x2 1 432 0 444 448 556 a3_x2
xsubckt_766_nand2_x0 1 0 1508 1525 1852 nand2_x0
xsubckt_818_nor2_x0 1 0 1462 1463 1466 nor2_x0
xsubckt_890_a4_x2 0 1402 1 1851 1854 1764 1762 a4_x2
xsubckt_606_a2_x2 0 77 1 78 425 a2_x2
xsubckt_147_a2_x2 0 529 1 530 546 a2_x2
xsubckt_137_a2_x2 0 539 1 542 548 a2_x2
xsubckt_688_ao22_x2 0 1581 1 646 47 1582 ao22_x2
xsubckt_408_nand2_x0 1 0 268 269 556 nand2_x0
xsubckt_1139_nand2_x0 1 0 1228 1229 239 nand2_x0
xsubckt_976_nand2_x0 1 0 1356 438 1757 nand2_x0
xsubckt_1871_sff1_x4 1 9 0 1613 1769 sff1_x4
xsubckt_1832_sff1_x4 1 9 0 1651 1794 sff1_x4
xsubckt_1401_a3_x2 1 1001 0 1002 1011 1020 a3_x2
xsubckt_1390_nand2_x0 1 0 1011 1013 1018 nand2_x0
xsubckt_1353_a4_x2 0 1045 1 1046 1047 1048 343 a4_x2
xsubckt_145_o2_x2 0 531 1 1800 1786 o2_x2
xsubckt_138_nand2_x0 1 0 538 542 548 nand2_x0
xsubckt_872_nand4_x0 1 0 1418 551 552 554 660 nand4_x0
xsubckt_940_mx2_x2 0 1696 1 1374 1830 1376 mx2_x2
xsubckt_1000_a2_x2 0 1336 1 412 505 a2_x2
xsubckt_1010_a2_x2 0 1326 1 1351 412 a2_x2
xsubckt_1471_a3_x2 1 934 0 935 79 369 a3_x2
xsubckt_1441_a3_x2 1 964 0 966 967 968 a3_x2
xsubckt_1349_nand2_x0 1 0 1049 1130 1767 nand2_x0
xsubckt_301_nand2_x0 1 0 375 383 495 nand2_x0
xsubckt_662_oa22_x2 0 23 1 281 360 631 oa22_x2
xsubckt_942_mx2_x2 0 1695 1 1373 1829 1412 mx2_x2
xsubckt_943_mx2_x2 0 1694 1 1373 1828 1403 mx2_x2
xsubckt_944_mx2_x2 0 1693 1 1373 1827 1398 mx2_x2
xsubckt_945_mx2_x2 0 1692 1 1373 1826 1394 mx2_x2
xsubckt_946_mx2_x2 0 1691 1 1373 1825 1393 mx2_x2
xsubckt_947_mx2_x2 0 1690 1 1373 1824 1385 mx2_x2
xsubckt_1273_ao22_x2 0 1117 1 651 1136 1118 ao22_x2
xsubckt_1867_sff1_x4 1 9 0 1617 1773 sff1_x4
xsubckt_1828_sff1_x4 1 9 0 1797 1805 sff1_x4
xsubckt_1718_ao22_x2 0 688 1 691 692 820 ao22_x2
xsubckt_1690_nand2_x0 1 0 716 718 963 nand2_x0
xsubckt_1344_a2_x2 0 1053 1 1054 1060 a2_x2
xsubckt_441_nor4_x0 1 0 236 237 238 242 461 nor4_x0
xsubckt_438_nand2_x0 1 0 239 473 495 nand2_x0
xsubckt_948_mx2_x2 0 1689 1 1373 1823 1380 mx2_x2
xsubckt_949_mx2_x2 0 1688 1 1373 1822 1376 mx2_x2
xsubckt_1032_nand2_x0 1 0 1669 1311 1313 nand2_x0
xsubckt_1159_a2_x2 0 1211 1 1212 1219 a2_x2
xsubckt_1658_a2_x2 0 748 1 749 925 a2_x2
xsubckt_1626_ao22_x2 0 780 1 784 786 940 ao22_x2
xsubckt_121_nand2_x0 1 0 555 655 1721 nand2_x0
xsubckt_992_nand4_x0 1 0 1344 420 504 517 520 nand4_x0
xsubckt_1056_mx2_x2 0 1662 1 438 1292 1747 mx2_x2
xsubckt_1189_a2_x2 0 1184 1 336 456 a2_x2
xsubckt_1775_sff1_x4 1 9 0 1699 1833 sff1_x4
xsubckt_1418_nand3_x0 1 0 986 545 550 1866 nand3_x0
xsubckt_1328_nand3_x0 1 0 1068 545 550 1858 nand3_x0
xsubckt_1379_nand2_x0 1 0 1021 1023 1028 nand2_x0
xsubckt_50_inv_x0 1 0 1780 618 inv_x0
xsubckt_51_inv_x0 1 0 1779 617 inv_x0
xsubckt_52_inv_x0 1 0 1874 616 inv_x0
xsubckt_53_inv_x0 1 0 1778 615 inv_x0
xsubckt_1192_nor4_x0 1 0 1181 1185 1187 1191 1192 nor4_x0
xsubckt_1646_o2_x2 0 760 1 762 764 o2_x2
xsubckt_454_nand4_x0 1 0 223 516 521 526 532 nand4_x0
xsubckt_54_inv_x0 1 0 1777 614 inv_x0
xsubckt_55_inv_x0 1 0 1776 613 inv_x0
xsubckt_56_inv_x0 1 0 1775 612 inv_x0
xsubckt_57_inv_x0 1 0 1865 611 inv_x0
xsubckt_58_inv_x0 1 0 1864 610 inv_x0
xsubckt_59_inv_x0 1 0 1863 609 inv_x0
xsubckt_318_a4_x2 0 358 1 588 1727 590 1729 a4_x2
xsubckt_919_nxr2_x1 1378 1 0 1390 642 nxr2_x1
xsubckt_985_nand3_x0 1 0 1349 1351 1365 413 nand3_x0
xsubckt_1062_nand2_x0 1 0 1660 1288 1290 nand2_x0
xsubckt_1185_nand4_x0 1 0 1188 551 586 1725 1728 nand4_x0
xsubckt_1674_nxr2_x1 732 1 0 733 915 nxr2_x1
xsubckt_1589_nand2_x0 1 0 817 819 1025 nand2_x0
xsubckt_1538_nand3_x0 1 0 868 481 554 1771 nand3_x0
xsubckt_426_a3_x2 1 251 0 415 417 420 a3_x2
xsubckt_200_a2_x2 0 476 1 1730 1729 a2_x2
xsubckt_717_nand3_x0 1 0 1555 58 63 1822 nand3_x0
xsubckt_1204_oa22_x2 0 1169 1 291 480 553 oa22_x2
xsubckt_1635_nxr2_x1 771 1 0 782 915 nxr2_x1
xsubckt_627_nand3_x0 1 0 56 57 64 1837 nand3_x0
xsubckt_524_a2_x2 0 154 1 155 156 a2_x2
xsubckt_329_a2_x2 0 347 1 348 350 a2_x2
xsubckt_905_a3_x2 1 1390 0 644 650 1762 a3_x2
xsubckt_1221_nand3_x0 1 0 1152 1155 74 334 nand3_x0
xsubckt_1278_oa22_x2 0 1113 1 1131 371 631 oa22_x2
xsubckt_785_nor2_x0 1 0 1491 1492 1495 nor2_x0
xsubckt_841_nand2_x0 1 0 1443 1458 1870 nand2_x0
xsubckt_1217_nand4_x0 1 0 1156 1157 1158 460 475 nand4_x0
xsubckt_1543_nxr2_x1 863 1 0 865 916 nxr2_x1
xsubckt_1431_nand3_x0 1 0 974 461 635 663 nand3_x0
xsubckt_498_nand2_x0 1 0 180 248 408 nand2_x0
xsubckt_216_nand4_x0 1 0 460 552 554 1730 591 nand4_x0
xsubckt_774_oa22_x2 0 1501 1 331 446 562 oa22_x2
xsubckt_978_nand2_x0 1 0 1677 1355 1356 nand2_x0
xsubckt_1891_sff1_x4 1 9 0 1593 1857 sff1_x4
xsubckt_1703_ao22_x2 0 703 1 705 707 765 ao22_x2
xsubckt_532_o2_x2 0 146 1 445 466 o2_x2
xsubckt_258_nor2_x0 1 0 418 1798 1786 nor2_x0
xsubckt_875_o4_x2 0 1415 1 1416 1417 73 355 o4_x2
xsubckt_1020_oa22_x2 0 1317 1 515 407 173 oa22_x2
xsubckt_1088_nand3_x0 1 0 1265 1266 1292 404 nand3_x0
xsubckt_1096_a4_x2 0 1258 1 1259 1260 1265 1334 a4_x2
xsubckt_1214_nand2_x0 1 0 1159 1160 491 nand2_x0
xsubckt_1852_sff1_x4 1 9 0 1632 1861 sff1_x4
xsubckt_1813_sff1_x4 1 9 0 1662 1747 sff1_x4
xsubckt_1438_a3_x2 1 967 0 1155 314 375 a3_x2
xsubckt_357_o2_x2 0 319 1 320 555 o2_x2
xsubckt_643_oa22_x2 0 1882 1 83 52 41 oa22_x2
xsubckt_657_nand3_x0 1 0 28 58 64 1843 nand3_x0
xsubckt_1037_a2_x2 0 1667 1 1306 1308 a2_x2
xsubckt_1887_sff1_x4 1 9 0 1597 1848 sff1_x4
xsubckt_1848_sff1_x4 1 9 0 1636 1865 sff1_x4
xsubckt_1809_sff1_x4 1 9 0 1666 1764 sff1_x4
xsubckt_1760_sff1_x4 1 9 0 1708 1818 sff1_x4
xsubckt_1701_a2_x2 0 705 1 768 772 a2_x2
xsubckt_1692_nand2_x0 1 0 714 722 731 nand2_x0
xsubckt_1282_a2_x2 0 1109 1 1110 1112 a2_x2
xsubckt_391_nand2_x0 1 0 285 286 290 nand2_x0
xsubckt_1034_nand2_x0 1 0 1308 438 657 nand2_x0
xsubckt_1057_a2_x2 0 1291 1 438 1723 a2_x2
xsubckt_1077_a2_x2 0 1658 1 1275 1284 a2_x2
xsubckt_1097_a2_x2 0 1257 1 1258 1271 a2_x2
xsubckt_1272_a2_x2 0 1118 1 1119 1120 a2_x2
xsubckt_603_nand2_x0 1 0 1720 80 83 nand2_x0
xsubckt_730_nand3_x0 1 0 1543 78 85 425 nand3_x0
xsubckt_1795_sff1_x4 1 9 0 1680 1737 sff1_x4
xsubckt_1756_sff1_x4 1 9 0 1712 1838 sff1_x4
xsubckt_1607_ao22_x2 0 799 1 912 802 905 ao22_x2
xsubckt_1596_a2_x2 0 810 1 811 812 a2_x2
xsubckt_1226_nor4_x0 1 0 1147 1148 1154 1156 1159 nor4_x0
xsubckt_1504_o2_x2 0 902 1 1855 1721 o2_x2
xsubckt_1281_nand3_x0 1 0 1110 1111 358 554 nand3_x0
xsubckt_421_a4_x2 0 256 1 413 419 504 538 a4_x2
xsubckt_419_nand3_x0 1 0 258 358 467 493 nand3_x0
xsubckt_333_nand2_x0 1 0 343 358 554 nand2_x0
xsubckt_687_nand3_x0 1 0 1582 358 547 554 nand3_x0
xsubckt_1197_ao22_x2 0 1176 1 495 493 338 ao22_x2
xsubckt_1712_oa22_x2 0 694 1 695 697 699 oa22_x2
xsubckt_1708_nxr2_x1 698 1 0 708 711 nxr2_x1
xsubckt_276_a4_x2 0 400 1 516 520 526 532 a4_x2
xsubckt_1031_ao22_x2 0 1309 1 533 527 439 ao22_x2
xsubckt_1064_nand2_x0 1 0 1286 1287 1342 nand2_x0
xsubckt_1491_nand3_x0 1 0 914 916 931 938 nand3_x0
xsubckt_153_nand2_x0 1 0 523 577 1786 nand2_x0
xsubckt_170_ao22_x2 0 506 1 1786 1796 546 ao22_x2
xsubckt_314_a3_x2 1 362 0 476 588 1727 a3_x2
xsubckt_670_nand3_x0 1 0 16 58 63 1826 nand3_x0
xsubckt_719_nand3_x0 1 0 1553 58 64 1838 nand3_x0
xsubckt_735_a4_x2 0 1538 1 551 586 1725 1727 a4_x2
xsubckt_755_a4_x2 0 1518 1 1519 1521 1522 1544 a4_x2
xsubckt_1224_oa22_x2 0 1149 1 1726 323 489 oa22_x2
xsubckt_629_nand3_x0 1 0 54 58 63 1829 nand3_x0
xsubckt_432_a2_x2 0 245 1 246 253 a2_x2
xsubckt_217_a2_x2 0 459 1 461 467 a2_x2
xsubckt_666_nand4_x0 1 0 19 20 21 22 23 nand4_x0
xsubckt_886_oa22_x2 0 1405 1 1408 1410 651 oa22_x2
xsubckt_1259_oa22_x2 0 1130 1 1133 1136 1144 oa22_x2
xsubckt_1497_ao22_x2 0 908 1 962 921 909 ao22_x2
xsubckt_1458_ao22_x2 0 947 1 642 953 949 ao22_x2
xsubckt_482_a2_x2 0 195 1 196 197 a2_x2
xsubckt_808_oa22_x2 0 1471 1 1521 1522 605 oa22_x2
xsubckt_843_nand2_x0 1 0 1441 1520 1850 nand2_x0
xsubckt_597_ao22_x2 0 85 1 494 337 279 ao22_x2
xsubckt_273_nand2_x0 1 0 403 516 520 nand2_x0
xsubckt_1039_nand4_x0 1 0 1304 551 554 1727 1721 nand4_x0
xsubckt_1128_nxr2_x1 1238 1 0 1846 1855 nxr2_x1
xsubckt_1443_a4_x2 0 962 1 964 969 973 978 a4_x2
xsubckt_1394_nand2_x0 1 0 1008 1137 1798 nand2_x0
xsubckt_1306_a3_x2 1 1087 0 1088 1097 1106 a3_x2
xsubckt_522_nand3_x0 1 0 156 362 493 556 nand3_x0
xsubckt_470_ao22_x2 0 207 1 215 211 208 ao22_x2
xsubckt_716_oa22_x2 0 1876 1 83 1561 1556 oa22_x2
xsubckt_1042_a3_x2 1 1301 0 1305 516 521 a3_x2
xsubckt_1872_sff1_x4 1 9 0 1612 1768 sff1_x4
xsubckt_1833_sff1_x4 1 9 0 1650 1793 sff1_x4
xsubckt_1606_nand2_x0 1 0 800 803 911 nand2_x0
xsubckt_1598_oa22_x2 0 808 1 811 812 939 oa22_x2
xsubckt_519_o2_x2 0 159 1 464 466 o2_x2
xsubckt_483_nand2_x0 1 0 194 196 197 nand2_x0
xsubckt_659_nand3_x0 1 0 26 58 63 1827 nand3_x0
xsubckt_951_mx2_x2 0 1687 1 1783 1372 345 mx2_x2
xsubckt_952_mx2_x2 0 1686 1 656 413 1754 mx2_x2
xsubckt_953_mx2_x2 0 1685 1 656 420 1753 mx2_x2
xsubckt_954_mx2_x2 0 1684 1 656 505 1752 mx2_x2
xsubckt_1110_a2_x2 0 1653 1 1247 1256 a2_x2
xsubckt_1126_nand2_x0 1 0 1240 1241 1242 nand2_x0
xsubckt_1868_sff1_x4 1 9 0 1616 1772 sff1_x4
xsubckt_1581_a3_x2 1 825 0 834 836 916 a3_x2
xsubckt_1571_a3_x2 1 835 0 932 937 1799 a3_x2
xsubckt_1434_a2_x2 0 971 1 1749 663 a2_x2
xsubckt_1432_oa22_x2 0 973 1 974 976 638 oa22_x2
xsubckt_1404_a2_x2 0 998 1 999 1000 a2_x2
xsubckt_479_nand3_x0 1 0 198 200 437 539 nand3_x0
xsubckt_186_nor2_x0 1 0 490 1728 1727 nor2_x0
xsubckt_1060_mx2_x2 0 1289 1 520 516 533 mx2_x2
xsubckt_1209_a2_x2 0 1164 1 79 331 a2_x2
xsubckt_1829_sff1_x4 1 9 0 1796 1804 sff1_x4
xsubckt_1780_sff1_x4 1 9 0 1694 1828 sff1_x4
xsubckt_1484_a2_x2 0 921 1 922 977 a2_x2
xsubckt_136_oa22_x2 0 540 1 667 560 545 oa22_x2
xsubckt_1066_mx2_x2 0 1659 1 438 1285 1748 mx2_x2
xsubckt_1776_sff1_x4 1 9 0 1698 1832 sff1_x4
xsubckt_1428_oa22_x2 0 977 1 1524 460 601 oa22_x2
xsubckt_1373_nand3_x0 1 0 1027 545 550 1870 nand3_x0
xsubckt_411_nand4_x0 1 0 265 275 554 655 1721 nand4_x0
xsubckt_1143_ao22_x2 0 1224 1 1225 1227 345 ao22_x2
xsubckt_1246_nand2_x0 1 0 1143 546 550 nand2_x0
xsubckt_548_nand4_x0 1 0 131 447 554 655 1721 nand4_x0
xsubckt_462_nand3_x0 1 0 215 481 554 556 nand3_x0
xsubckt_60_inv_x0 1 0 1862 608 inv_x0
xsubckt_243_ao22_x2 0 433 1 513 502 435 ao22_x2
xsubckt_993_nand2_x0 1 0 1343 1344 1347 nand2_x0
xsubckt_1105_nand3_x0 1 0 1251 173 411 525 nand3_x0
xsubckt_1732_oa22_x2 0 674 1 675 678 656 oa22_x2
xsubckt_1728_nxr2_x1 678 1 0 679 682 nxr2_x1
xsubckt_1574_ao22_x2 0 832 1 835 837 940 ao22_x2
xsubckt_1294_nor2_x0 1 0 1098 1099 1102 nor2_x0
xsubckt_440_oa22_x2 0 237 1 495 292 387 oa22_x2
xsubckt_61_inv_x0 1 0 1861 607 inv_x0
xsubckt_62_inv_x0 1 0 1860 606 inv_x0
xsubckt_63_inv_x0 1 0 1859 605 inv_x0
xsubckt_64_inv_x0 1 0 1858 604 inv_x0
xsubckt_65_inv_x0 1 0 1746 603 inv_x0
xsubckt_66_inv_x0 1 0 1784 602 inv_x0
xsubckt_174_a4_x2 0 502 1 505 520 526 532 a4_x2
xsubckt_231_nand4_x0 1 0 445 551 554 1728 589 nand4_x0
xsubckt_852_nand3_x0 1 0 1434 1518 1526 1777 nand3_x0
xsubckt_1746_o2_x2 0 669 1 692 656 o2_x2
xsubckt_1442_nand4_x0 1 0 963 965 967 969 973 nand4_x0
xsubckt_621_nand4_x0 1 0 62 551 552 554 1751 nand4_x0
xsubckt_67_inv_x0 1 0 1733 601 inv_x0
xsubckt_68_inv_x0 1 0 1804 600 inv_x0
xsubckt_69_inv_x0 1 0 1883 599 inv_x0
xsubckt_192_nand3_x0 1 0 484 552 590 1729 nand3_x0
xsubckt_232_a3_x2 1 444 0 445 446 452 a3_x2
xsubckt_252_a3_x2 1 424 0 467 481 495 a3_x2
xsubckt_278_nand4_x0 1 0 398 402 404 405 437 nand4_x0
xsubckt_1640_oa22_x2 0 766 1 911 771 906 oa22_x2
xsubckt_1636_nxr2_x1 770 1 0 782 916 nxr2_x1
xsubckt_1366_nand2_x0 1 0 1033 1034 1040 nand2_x0
xsubckt_566_a3_x2 1 113 0 114 118 119 a3_x2
xsubckt_536_a3_x2 1 142 0 143 148 149 a3_x2
xsubckt_526_a3_x2 1 152 0 154 157 161 a3_x2
xsubckt_155_a2_x2 0 521 1 522 523 a2_x2
xsubckt_469_a2_x2 0 208 1 209 210 a2_x2
xsubckt_845_nand2_x0 1 0 1903 1440 1444 nand2_x0
xsubckt_1198_nor2_x0 1 0 1175 1176 321 nor2_x0
xsubckt_1312_ao22_x2 0 1082 1 645 1136 1084 ao22_x2
xsubckt_250_o3_x2 0 426 1 428 433 440 o3_x2
xsubckt_275_nand2_x0 1 0 401 526 532 nand2_x0
xsubckt_747_nor2_x0 1 0 1526 1527 1535 nor2_x0
xsubckt_1136_a4_x2 0 1231 1 473 495 585 641 a4_x2
xsubckt_534_o3_x2 0 144 1 145 474 555 o3_x2
xsubckt_123_o2_x2 0 553 1 1726 1725 o2_x2
xsubckt_1186_a4_x2 0 1187 1 551 586 1725 1728 a4_x2
xsubckt_1853_sff1_x4 1 9 0 1631 1860 sff1_x4
xsubckt_1814_sff1_x4 1 9 0 1661 1723 sff1_x4
xsubckt_1518_a3_x2 1 888 0 889 890 911 a3_x2
xsubckt_248_oa22_x2 0 428 1 477 432 429 oa22_x2
xsubckt_307_nand2_x0 1 0 369 383 554 nand2_x0
xsubckt_1888_sff1_x4 1 9 0 1596 1847 sff1_x4
xsubckt_1308_mx2_x2 0 1616 1 656 1086 1772 mx2_x2
xsubckt_395_nand2_x0 1 0 281 292 554 nand2_x0
xsubckt_965_nand2_x0 1 0 1681 1364 1366 nand2_x0
xsubckt_1255_ao22_x2 0 1134 1 553 357 371 ao22_x2
xsubckt_1849_sff1_x4 1 9 0 1635 1864 sff1_x4
xsubckt_1761_sff1_x4 1 9 0 1707 1817 sff1_x4
xsubckt_1657_mx2_x2 0 749 1 752 927 940 mx2_x2
xsubckt_607_nand2_x0 1 0 76 78 425 nand2_x0
xsubckt_644_nand3_x0 1 0 40 57 63 1820 nand3_x0
xsubckt_679_oa22_x2 0 1879 1 83 13 1590 oa22_x2
xsubckt_1187_a2_x2 0 1186 1 274 287 a2_x2
xsubckt_1201_nand2_x0 1 0 1172 68 85 nand2_x0
xsubckt_1796_sff1_x4 1 9 0 1679 1758 sff1_x4
xsubckt_1696_a2_x2 0 710 1 741 743 a2_x2
xsubckt_1647_ao22_x2 0 759 1 36 957 761 ao22_x2
xsubckt_1375_nand3_x0 1 0 1025 383 554 1870 nand3_x0
xsubckt_1338_nand2_x0 1 0 1059 1137 1803 nand2_x0
xsubckt_554_nand3_x0 1 0 125 275 467 554 nand3_x0
xsubckt_517_nand2_x0 1 0 161 211 216 nand2_x0
xsubckt_1021_nand2_x0 1 0 1316 1317 504 nand2_x0
xsubckt_1127_xr2_x1 1239 0 1 1857 1856 xr2_x1
xsubckt_1268_mx2_x2 0 1620 1 656 1122 1782 mx2_x2
xsubckt_1757_sff1_x4 1 9 0 1711 1821 sff1_x4
xsubckt_1638_nand2_x0 1 0 768 771 911 nand2_x0
xsubckt_1501_nand2_x0 1 0 904 905 909 nand2_x0
xsubckt_1317_nxr2_x1 1077 1 0 1080 1087 nxr2_x1
xsubckt_1107_nand3_x0 1 0 1249 1250 503 527 nand3_x0
xsubckt_1614_o2_x2 0 792 1 951 562 o2_x2
xsubckt_1555_ao22_x2 0 851 1 867 869 940 ao22_x2
xsubckt_1321_nand2_x0 1 0 1074 1076 343 nand2_x0
xsubckt_247_nand2_x0 1 0 429 430 454 nand2_x0
xsubckt_817_nand2_x0 1 0 1463 1464 1465 nand2_x0
xsubckt_1709_nxr2_x1 697 1 0 708 712 nxr2_x1
xsubckt_1444_nand4_x0 1 0 961 964 969 973 978 nand4_x0
xsubckt_1407_nand3_x0 1 0 996 545 550 1867 nand3_x0
xsubckt_410_nand2_x0 1 0 266 275 554 nand2_x0
xsubckt_366_a4_x2 0 310 1 476 490 586 1725 a4_x2
xsubckt_157_nand2_x0 1 0 519 574 1786 nand2_x0
xsubckt_1264_oa22_x2 0 1125 1 1853 1135 1126 oa22_x2
xsubckt_584_nand3_x0 1 0 4 97 104 228 nand3_x0
xsubckt_502_a2_x2 0 176 1 177 255 a2_x2
xsubckt_494_a3_x2 1 184 0 223 226 295 a3_x2
xsubckt_457_nand2_x0 1 0 220 310 556 nand2_x0
xsubckt_327_a2_x2 0 349 1 358 495 a2_x2
xsubckt_320_nand2_x0 1 0 356 358 587 nand2_x0
xsubckt_887_nxr2_x1 1404 1 0 1407 1852 nxr2_x1
xsubckt_903_a3_x2 1 1392 0 1855 1764 1762 a3_x2
xsubckt_923_a3_x2 1 1375 0 1414 57 63 a3_x2
xsubckt_1028_ao22_x2 0 1312 1 511 507 439 ao22_x2
xsubckt_1695_oa22_x2 0 711 1 714 717 721 oa22_x2
xsubckt_1668_nand2_x0 1 0 738 740 744 nand2_x0
xsubckt_1656_oa22_x2 0 750 1 754 756 939 oa22_x2
xsubckt_1531_nand2_x0 1 0 875 876 877 nand2_x0
xsubckt_562_a2_x2 0 117 1 118 119 a2_x2
xsubckt_140_nand2_x0 1 0 536 571 1786 nand2_x0
xsubckt_974_nand3_x0 1 0 1357 1360 1365 413 nand3_x0
xsubckt_983_a3_x2 1 1351 0 419 506 509 a3_x2
xsubckt_1188_nand2_x0 1 0 1185 274 287 nand2_x0
xsubckt_1351_nand2_x0 1 0 1047 372 1852 nand2_x0
xsubckt_620_nand2_x0 1 0 63 66 70 nand2_x0
xsubckt_706_nand3_x0 1 0 1565 58 64 1839 nand3_x0
xsubckt_809_oa22_x2 0 1470 1 331 446 558 oa22_x2
xsubckt_847_nand2_x0 1 0 1438 1458 1869 nand2_x0
xsubckt_1129_nxr2_x1 1237 1 0 1238 1239 nxr2_x1
xsubckt_876_a2_x2 0 1414 1 1415 1721 a2_x2
xsubckt_1261_nand2_x0 1 0 1128 1131 371 nand2_x0
xsubckt_1873_sff1_x4 1 9 0 1611 1767 sff1_x4
xsubckt_1724_ao22_x2 0 682 1 684 685 870 ao22_x2
xsubckt_1398_a4_x2 0 1004 1 1005 1006 1007 343 a4_x2
xsubckt_260_nand2_x0 1 0 416 592 1786 nand2_x0
xsubckt_804_o2_x2 0 1895 1 1475 1482 o2_x2
xsubckt_830_nand2_x0 1 0 1452 1531 1802 nand2_x0
xsubckt_960_mx2_x2 0 1367 1 438 419 1741 mx2_x2
xsubckt_1834_sff1_x4 1 9 0 1649 1792 sff1_x4
xsubckt_1671_a3_x2 1 735 0 932 937 1803 a3_x2
xsubckt_1651_a3_x2 1 755 0 932 937 1802 a3_x2
xsubckt_1420_nand3_x0 1 0 984 383 554 1866 nand3_x0
xsubckt_346_nand3_x0 1 0 330 338 493 556 nand3_x0
xsubckt_664_oa22_x2 0 21 1 48 482 648 oa22_x2
xsubckt_874_o2_x2 0 1416 1 1538 457 o2_x2
xsubckt_1012_o4_x2 0 1324 1 1327 1333 1339 1343 o4_x2
xsubckt_1055_a2_x2 0 1292 1 1351 413 a2_x2
xsubckt_1075_a2_x2 0 1276 1 1277 439 a2_x2
xsubckt_1115_mx2_x2 0 1651 1 1246 1803 1794 mx2_x2
xsubckt_1116_mx2_x2 0 1650 1 1246 1802 1793 mx2_x2
xsubckt_1260_a2_x2 0 1129 1 1131 371 a2_x2
xsubckt_1869_sff1_x4 1 9 0 1615 1771 sff1_x4
xsubckt_1781_sff1_x4 1 9 0 1693 1827 sff1_x4
xsubckt_1564_a2_x2 0 842 1 853 978 a2_x2
xsubckt_1557_nand3_x0 1 0 849 866 868 927 nand3_x0
xsubckt_1544_a2_x2 0 862 1 864 911 a2_x2
xsubckt_1524_a2_x2 0 882 1 883 884 a2_x2
xsubckt_1467_nand3_x0 1 0 938 481 554 1769 nand3_x0
xsubckt_176_oa22_x2 0 500 1 501 512 539 oa22_x2
xsubckt_1085_a2_x2 0 1657 1 1268 1274 a2_x2
xsubckt_1117_mx2_x2 0 1649 1 1246 1801 1792 mx2_x2
xsubckt_1118_mx2_x2 0 1648 1 1246 1800 1791 mx2_x2
xsubckt_1119_mx2_x2 0 1647 1 1246 1799 1790 mx2_x2
xsubckt_1429_oa22_x2 0 976 1 1524 460 634 oa22_x2
xsubckt_1399_a2_x2 0 1003 1 1004 1008 a2_x2
xsubckt_1389_a2_x2 0 1012 1 1013 1018 a2_x2
xsubckt_646_nand3_x0 1 0 38 58 64 1844 nand3_x0
xsubckt_1113_nand2_x0 1 0 1244 1245 438 nand2_x0
xsubckt_1150_nand3_x0 1 0 1219 377 482 549 nand3_x0
xsubckt_1777_sff1_x4 1 9 0 1697 1831 sff1_x4
xsubckt_1540_nand3_x0 1 0 866 932 937 1798 nand3_x0
xsubckt_593_nand4_x0 1 0 88 383 467 586 1725 nand4_x0
xsubckt_860_nand2_x0 1 0 1427 1531 1797 nand2_x0
xsubckt_1413_nand2_x0 1 0 990 992 997 nand2_x0
xsubckt_529_oa22_x2 0 149 1 166 167 436 oa22_x2
xsubckt_70_inv_x0 1 0 1787 598 inv_x0
xsubckt_71_inv_x0 1 0 1805 597 inv_x0
xsubckt_72_inv_x0 1 0 1884 596 inv_x0
xsubckt_73_inv_x0 1 0 1788 595 inv_x0
xsubckt_205_ao22_x2 0 471 1 492 472 474 ao22_x2
xsubckt_715_nand4_x0 1 0 1556 1557 1558 1559 1560 nand4_x0
xsubckt_819_nand2_x0 1 0 1461 1462 1467 nand2_x0
xsubckt_1729_nxr2_x1 677 1 0 686 688 nxr2_x1
xsubckt_1409_nand3_x0 1 0 994 383 554 1867 nand3_x0
xsubckt_1319_nand3_x0 1 0 1076 545 550 1859 nand3_x0
xsubckt_568_a4_x2 0 111 1 112 205 260 390 a4_x2
xsubckt_558_a4_x2 0 121 1 122 189 198 201 a4_x2
xsubckt_74_inv_x0 1 0 1806 594 inv_x0
xsubckt_75_inv_x0 1 0 1885 593 inv_x0
xsubckt_76_inv_x0 1 0 1789 592 inv_x0
xsubckt_77_inv_x0 1 0 1729 591 inv_x0
xsubckt_78_inv_x0 1 0 1730 590 inv_x0
xsubckt_79_inv_x0 1 0 1727 589 inv_x0
xsubckt_1270_nand3_x0 1 0 1120 545 550 1864 nand3_x0
xsubckt_578_a4_x2 0 102 1 353 359 394 395 a4_x2
xsubckt_322_nand2_x0 1 0 354 358 493 nand2_x0
xsubckt_177_a3_x2 1 499 0 552 1730 591 a3_x2
xsubckt_187_a3_x2 1 489 0 490 1730 591 a3_x2
xsubckt_225_a2_x2 0 451 1 1726 1725 a2_x2
xsubckt_811_a3_x2 1 1468 0 1469 1472 1473 a3_x2
xsubckt_1002_nand3_x0 1 0 1334 1336 1338 525 nand3_x0
xsubckt_1053_nand2_x0 1 0 1293 1294 1295 nand2_x0
xsubckt_1676_oa22_x2 0 730 1 911 732 906 oa22_x2
xsubckt_1570_nand3_x0 1 0 836 481 554 1772 nand3_x0
xsubckt_460_a2_x2 0 217 1 218 222 a2_x2
xsubckt_369_nand2_x0 1 0 307 310 467 nand2_x0
xsubckt_148_ao22_x2 0 528 1 1786 1800 546 ao22_x2
xsubckt_265_a2_x2 0 411 1 504 538 a2_x2
xsubckt_1480_nand3_x0 1 0 925 928 941 943 nand3_x0
xsubckt_579_a2_x2 0 101 1 102 103 a2_x2
xsubckt_549_a2_x2 0 130 1 131 132 a2_x2
xsubckt_702_oa22_x2 0 1568 1 281 360 628 oa22_x2
xsubckt_708_nand3_x0 1 0 1563 58 63 1823 nand3_x0
xsubckt_744_a2_x2 0 1529 1 325 334 a2_x2
xsubckt_849_nand2_x0 1 0 1436 1520 1849 nand2_x0
xsubckt_1421_a4_x2 0 983 1 984 985 986 343 a4_x2
xsubckt_390_o3_x2 0 286 1 287 555 587 o3_x2
xsubckt_175_nand4_x0 1 0 501 505 520 526 532 nand4_x0
xsubckt_213_o2_x2 0 463 1 464 555 o2_x2
xsubckt_1030_a3_x2 1 1310 0 504 517 520 a3_x2
xsubckt_1702_mx2_x2 0 704 1 772 767 769 mx2_x2
xsubckt_1296_a4_x2 0 1096 1 1097 1107 1115 1124 a4_x2
xsubckt_537_o2_x2 0 141 1 334 555 o2_x2
xsubckt_211_nand3_x0 1 0 465 467 497 1725 nand3_x0
xsubckt_1090_a3_x2 1 1263 0 1264 1265 1334 a3_x2
xsubckt_1854_sff1_x4 1 9 0 1630 1859 sff1_x4
xsubckt_1815_sff1_x4 1 9 0 1660 1724 sff1_x4
xsubckt_1563_nand2_x0 1 0 843 845 859 nand2_x0
xsubckt_1492_oa22_x2 0 913 1 938 931 916 oa22_x2
xsubckt_1412_a2_x2 0 991 1 992 997 a2_x2
xsubckt_601_nand3_x0 1 0 81 444 479 487 nand3_x0
xsubckt_475_nand4_x0 1 0 202 402 437 515 539 nand4_x0
xsubckt_385_nand4_x0 1 0 291 588 1727 1730 591 nand4_x0
xsubckt_172_nand2_x0 1 0 504 508 510 nand2_x0
xsubckt_262_nand2_x0 1 0 414 416 546 nand2_x0
xsubckt_828_nand3_x0 1 0 1454 1518 1526 1767 nand3_x0
xsubckt_969_nand2_x0 1 0 1361 438 1758 nand2_x0
xsubckt_1079_nand3_x0 1 0 1273 1326 173 401 nand3_x0
xsubckt_1199_a3_x2 1 1174 0 1175 1177 1179 a3_x2
xsubckt_1889_sff1_x4 1 9 0 1595 1846 sff1_x4
xsubckt_1762_sff1_x4 1 9 0 1706 1816 sff1_x4
xsubckt_1706_a2_x2 0 700 1 461 1764 a2_x2
xsubckt_1663_mx2_x2 0 743 1 978 746 788 mx2_x2
xsubckt_1662_mx2_x2 0 744 1 978 745 787 mx2_x2
xsubckt_1661_mx2_x2 0 745 1 759 747 751 mx2_x2
xsubckt_1660_mx2_x2 0 746 1 759 748 750 mx2_x2
xsubckt_1613_ao22_x2 0 793 1 954 1540 1851 ao22_x2
xsubckt_1482_a2_x2 0 923 1 924 925 a2_x2
xsubckt_1472_a2_x2 0 933 1 1158 1189 a2_x2
xsubckt_1452_a2_x2 0 953 1 955 1541 a2_x2
xsubckt_1383_nand2_x0 1 0 1018 1130 1778 nand2_x0
xsubckt_1318_mx2_x2 0 1615 1 656 1077 1771 mx2_x2
xsubckt_129_nor2_x0 1 0 547 1874 1783 nor2_x0
xsubckt_738_nand3_x0 1 0 1535 1537 1539 1541 nand3_x0
xsubckt_1687_ao22_x2 0 719 1 918 917 912 ao22_x2
xsubckt_599_nor2_x0 1 0 83 84 483 nor2_x0
xsubckt_685_nand4_x0 1 0 1584 1586 1587 1588 1589 nand4_x0
xsubckt_1277_mx2_x2 0 1619 1 656 1114 1781 mx2_x2
xsubckt_1797_sff1_x4 1 9 0 1678 1736 sff1_x4
xsubckt_1758_sff1_x4 1 9 0 1710 1820 sff1_x4
xsubckt_1357_nxr2_x1 1041 1 0 1043 1051 nxr2_x1
xsubckt_468_nand3_x0 1 0 209 383 467 586 nand3_x0
xsubckt_417_nand4_x0 1 0 259 261 293 304 311 nand4_x0
xsubckt_1679_nand3_x0 1 0 727 734 736 927 nand3_x0
xsubckt_1295_o2_x2 0 1097 1 1099 1102 o2_x2
xsubckt_611_a4_x2 0 72 1 316 345 456 464 a4_x2
xsubckt_416_a4_x2 0 260 1 261 293 304 311 a4_x2
xsubckt_858_nand3_x0 1 0 1429 1518 1526 1776 nand3_x0
xsubckt_999_nand2_x0 1 0 1337 1338 525 nand2_x0
xsubckt_1362_nand3_x0 1 0 1037 383 554 1871 nand3_x0
xsubckt_504_nand2_x0 1 0 174 175 232 nand2_x0
xsubckt_288_nand3_x0 1 0 388 476 1728 589 nand3_x0
xsubckt_892_nxr2_x1 1400 1 0 1411 648 nxr2_x1
xsubckt_1625_nand2_x0 1 0 781 783 785 nand2_x0
xsubckt_514_a3_x2 1 164 0 165 199 230 a3_x2
xsubckt_451_nand3_x0 1 0 226 257 404 525 nand3_x0
xsubckt_359_a3_x2 1 317 0 447 1726 587 a3_x2
xsubckt_143_a2_x2 0 533 1 535 537 a2_x2
xsubckt_982_nand2_x0 1 0 1352 438 1756 nand2_x0
xsubckt_1572_nand3_x0 1 0 834 932 937 1799 nand3_x0
xsubckt_594_a3_x2 1 87 0 88 89 126 a3_x2
xsubckt_437_a2_x2 0 240 1 473 495 a2_x2
xsubckt_144_nand2_x0 1 0 532 535 537 nand2_x0
xsubckt_183_a2_x2 0 493 1 1726 587 a2_x2
xsubckt_193_a2_x2 0 483 1 485 495 a2_x2
xsubckt_220_nand4_x0 1 0 456 551 552 1726 587 nand4_x0
xsubckt_838_a3_x2 1 1445 0 1446 1447 1448 a3_x2
xsubckt_520_nand4_x0 1 0 158 467 551 552 554 nand4_x0
xsubckt_868_a3_x2 1 1420 0 1421 1422 1423 a3_x2
xsubckt_1745_nand2_x0 1 0 670 1854 656 nand2_x0
xsubckt_430_nand4_x0 1 0 247 249 402 404 437 nand4_x0
xsubckt_206_nor2_x0 1 0 470 1724 1855 nor2_x0
xsubckt_1124_nand3_x0 1 0 1242 1243 377 549 nand3_x0
xsubckt_1800_sff1_x4 1 9 0 1675 1756 sff1_x4
xsubckt_1468_a4_x2 0 937 1 1155 1169 314 375 a4_x2
xsubckt_625_mx2_x2 0 58 1 65 60 584 mx2_x2
xsubckt_481_nand3_x0 1 0 196 358 467 554 nand3_x0
xsubckt_340_nand4_x0 1 0 336 490 554 590 1729 nand4_x0
xsubckt_956_ao22_x2 0 1370 1 545 422 439 ao22_x2
xsubckt_1874_sff1_x4 1 9 0 1610 1780 sff1_x4
xsubckt_1835_sff1_x4 1 9 0 1648 1791 sff1_x4
xsubckt_1565_nand2_x0 1 0 841 853 978 nand2_x0
xsubckt_1320_a2_x2 0 1075 1 1076 343 a2_x2
xsubckt_1310_a2_x2 0 1084 1 1085 343 a2_x2
xsubckt_1300_a2_x2 0 1093 1 1094 343 a2_x2
xsubckt_626_mx2_x2 0 57 1 65 59 1732 mx2_x2
xsubckt_264_nand2_x0 1 0 412 415 417 nand2_x0
xsubckt_650_o2_x2 0 34 1 51 619 o2_x2
xsubckt_665_oa22_x2 0 20 1 44 343 668 oa22_x2
xsubckt_957_nand4_x0 1 0 1369 1370 257 404 525 nand4_x0
xsubckt_1120_mx2_x2 0 1646 1 1246 1798 1789 mx2_x2
xsubckt_1121_mx2_x2 0 1645 1 1246 1797 1788 mx2_x2
xsubckt_1122_mx2_x2 0 1644 1 1246 1796 1787 mx2_x2
xsubckt_1624_a2_x2 0 782 1 783 785 a2_x2
xsubckt_1475_nand2_x0 1 0 930 931 938 nand2_x0
xsubckt_1381_nxr2_x1 1019 1 0 1022 1032 nxr2_x1
xsubckt_1370_a2_x2 0 1029 1 1030 1031 a2_x2
xsubckt_825_ao22_x2 0 1456 1 652 1521 1544 ao22_x2
xsubckt_1195_a2_x2 0 1178 1 381 482 a2_x2
xsubckt_1782_sff1_x4 1 9 0 1692 1826 sff1_x4
xsubckt_1469_a2_x2 0 936 1 85 302 a2_x2
xsubckt_423_nand3_x0 1 0 254 256 402 404 nand3_x0
xsubckt_1184_ao22_x2 0 1189 1 494 472 456 ao22_x2
xsubckt_1778_sff1_x4 1 9 0 1696 1830 sff1_x4
xsubckt_1507_nand2_x0 1 0 899 900 1057 nand2_x0
xsubckt_1303_oa22_x2 0 1090 1 1849 1135 1092 oa22_x2
xsubckt_813_nand3_x0 1 0 1467 1518 1526 1769 nand3_x0
xsubckt_1013_nand4_x0 1 0 1323 250 504 516 521 nand4_x0
xsubckt_1027_nand2_x0 1 0 1313 438 1738 nand2_x0
xsubckt_1106_ao22_x2 0 1250 1 414 418 419 ao22_x2
xsubckt_1584_o3_x2 0 822 1 824 825 912 o3_x2
xsubckt_1502_ao22_x2 0 903 1 906 910 1721 ao22_x2
xsubckt_1447_o2_x2 0 958 1 960 975 o2_x2
xsubckt_1417_nand2_x0 1 0 987 1130 1775 nand2_x0
xsubckt_80_inv_x0 1 0 1728 588 inv_x0
xsubckt_304_a4_x2 0 372 1 476 554 1728 589 a4_x2
xsubckt_1734_oa22_x2 0 673 1 720 714 717 oa22_x2
xsubckt_618_a4_x2 0 65 1 67 71 77 549 a4_x2
xsubckt_384_a4_x2 0 292 1 588 1727 1730 591 a4_x2
xsubckt_86_inv_x0 1 0 1748 582 inv_x0
xsubckt_85_inv_x0 1 0 1751 583 inv_x0
xsubckt_84_inv_x0 1 0 1732 584 inv_x0
xsubckt_83_inv_x0 1 0 1735 585 inv_x0
xsubckt_82_inv_x0 1 0 1726 586 inv_x0
xsubckt_81_inv_x0 1 0 1725 587 inv_x0
xsubckt_179_a4_x2 0 497 1 552 586 1730 591 a4_x2
xsubckt_1100_nand2_x0 1 0 1256 438 603 nand2_x0
xsubckt_1603_nxr2_x1 803 1 0 810 915 nxr2_x1
xsubckt_1400_nand2_x0 1 0 1002 1003 1009 nand2_x0
xsubckt_500_a2_x2 0 178 1 179 500 a2_x2
xsubckt_472_a3_x2 1 205 0 206 228 245 a3_x2
xsubckt_363_nand3_x0 1 0 313 323 556 1726 nand3_x0
xsubckt_89_inv_x0 1 0 1811 579 inv_x0
xsubckt_88_inv_x0 1 0 1750 580 inv_x0
xsubckt_87_inv_x0 1 0 1731 581 inv_x0
xsubckt_267_a3_x2 1 409 0 412 504 538 a3_x2
xsubckt_277_a3_x2 1 399 0 402 404 405 a3_x2
xsubckt_287_a3_x2 1 389 0 476 1728 589 a3_x2
xsubckt_648_a4_x2 0 36 1 37 38 39 40 a4_x2
xsubckt_698_a4_x2 0 1572 1 1574 1575 1576 1577 a4_x2
xsubckt_1006_nand3_x0 1 0 1330 1360 412 538 nand3_x0
xsubckt_1133_nand4_x0 1 0 1233 1234 551 552 554 nand4_x0
xsubckt_1688_nor2_x0 1 0 718 719 978 nor2_x0
xsubckt_637_ao22_x2 0 46 1 338 485 495 ao22_x2
xsubckt_609_a2_x2 0 74 1 316 345 a2_x2
xsubckt_550_a2_x2 0 129 1 130 133 a2_x2
xsubckt_736_a3_x2 1 1537 0 316 360 377 a3_x2
xsubckt_753_nand3_x0 1 0 1520 371 445 479 nand3_x0
xsubckt_941_a3_x2 1 1373 0 1414 58 63 a3_x2
xsubckt_619_a2_x2 0 64 1 66 70 a2_x2
xsubckt_570_a2_x2 0 109 1 110 340 a2_x2
xsubckt_146_nand2_x0 1 0 530 568 1786 nand2_x0
xsubckt_1747_nand2_x0 1 0 1594 669 670 nand2_x0
xsubckt_1316_a4_x2 0 1078 1 1079 1088 1097 1106 a4_x2
xsubckt_1314_ao22_x2 0 1080 1 628 1129 1082 ao22_x2
xsubckt_884_a2_x2 0 1407 1 1408 1410 a2_x2
xsubckt_1040_nand2_x0 1 0 1303 1304 1764 nand2_x0
xsubckt_1820_sff1_x4 1 9 0 1655 1750 sff1_x4
xsubckt_1388_ao22_x2 0 1013 1 560 1138 1014 ao22_x2
xsubckt_1376_a4_x2 0 1024 1 1025 1026 1027 343 a4_x2
xsubckt_1346_a4_x2 0 1051 1 1052 1065 1070 1078 a4_x2
xsubckt_393_nand3_x0 1 0 283 289 493 556 nand3_x0
xsubckt_343_o2_x2 0 333 1 334 466 o2_x2
xsubckt_342_nand4_x0 1 0 334 476 490 1726 587 nand4_x0
xsubckt_128_o2_x2 0 548 1 1799 1786 o2_x2
xsubckt_802_o2_x2 0 1476 1 1477 1480 o2_x2
xsubckt_836_nand2_x0 1 0 1447 1520 1851 nand2_x0
xsubckt_912_nand4_x0 1 0 1384 1847 1855 1764 1762 nand4_x0
xsubckt_1036_nand3_x0 1 0 1306 1307 1328 439 nand3_x0
xsubckt_1855_sff1_x4 1 9 0 1629 1858 sff1_x4
xsubckt_1816_sff1_x4 1 9 0 1659 1748 sff1_x4
xsubckt_1516_nand3_x0 1 0 890 891 893 916 nand3_x0
xsubckt_1439_nor3_x0 1 0 966 1161 332 349 nor3_x0
xsubckt_1415_nxr2_x1 988 1 0 991 1001 nxr2_x1
xsubckt_605_nand3_x0 1 0 78 358 450 553 nand3_x0
xsubckt_389_nand4_x0 1 0 287 551 586 588 1727 nand4_x0
xsubckt_266_nand2_x0 1 0 410 504 538 nand2_x0
xsubckt_1063_a2_x2 0 1287 1 1351 539 a2_x2
xsubckt_1087_nand2_x0 1 0 1266 532 539 nand2_x0
xsubckt_1249_a3_x2 1 1140 0 1141 297 336 a3_x2
xsubckt_1532_a2_x2 0 874 1 875 925 a2_x2
xsubckt_1327_mx2_x2 0 1614 1 656 1069 1770 mx2_x2
xsubckt_642_nand4_x0 1 0 41 42 45 49 50 nand4_x0
xsubckt_693_nand3_x0 1 0 1577 58 63 1824 nand3_x0
xsubckt_1058_oa22_x2 0 1661 1 1350 1295 1291 oa22_x2
xsubckt_1093_a2_x2 0 1261 1 438 580 a2_x2
xsubckt_1109_o4_x2 0 1247 1 1248 1252 1254 1270 o4_x2
xsubckt_1218_ao22_x2 0 1155 1 494 388 325 ao22_x2
xsubckt_1763_sff1_x4 1 9 0 1705 1815 sff1_x4
xsubckt_1550_nand2_x0 1 0 856 858 1006 nand2_x0
xsubckt_425_nand3_x0 1 0 252 358 467 495 nand3_x0
xsubckt_1798_sff1_x4 1 9 0 1677 1757 sff1_x4
xsubckt_1323_oa22_x2 0 1072 1 1847 1135 1074 oa22_x2
xsubckt_1289_mx2_x2 0 1618 1 656 1103 1774 mx2_x2
xsubckt_245_nand3_x0 1 0 431 470 655 1721 nand3_x0
xsubckt_866_nand2_x0 1 0 1422 1531 1796 nand2_x0
xsubckt_1015_nand4_x0 1 0 1321 412 504 516 521 nand4_x0
xsubckt_1759_sff1_x4 1 9 0 1709 1819 sff1_x4
xsubckt_1597_nand2_x0 1 0 809 811 812 nand2_x0
xsubckt_1419_nand2_x0 1 0 985 372 1846 nand2_x0
xsubckt_635_nand3_x0 1 0 48 338 495 621 nand3_x0
xsubckt_222_a4_x2 0 454 1 455 458 463 465 a4_x2
xsubckt_282_nand4_x0 1 0 394 469 473 493 556 nand4_x0
xsubckt_1609_o2_x2 0 797 1 799 804 o2_x2
xsubckt_1329_nand2_x0 1 0 1067 1068 343 nand2_x0
xsubckt_622_ao22_x2 0 61 1 582 67 62 ao22_x2
xsubckt_545_nand3_x0 1 0 134 275 451 467 nand3_x0
xsubckt_508_nand2_x0 1 0 170 171 172 nand2_x0
xsubckt_404_nand4_x0 1 0 272 275 451 655 1721 nand4_x0
xsubckt_310_a3_x2 1 366 0 368 655 1721 a3_x2
xsubckt_721_a4_x2 0 1551 1 1552 1553 1554 1555 a4_x2
xsubckt_741_a4_x2 0 1532 1 1534 385 453 471 a4_x2
xsubckt_749_ao22_x2 0 1524 1 494 472 309 ao22_x2
xsubckt_893_nxr2_x1 1399 1 0 1400 1405 nxr2_x1
xsubckt_1190_nand2_x0 1 0 1183 336 456 nand2_x0
xsubckt_1280_nand2_x0 1 0 1111 1783 666 nand2_x0
xsubckt_1580_nand2_x0 1 0 826 828 831 nand2_x0
xsubckt_586_a4_x2 0 95 1 247 252 298 301 a4_x2
xsubckt_986_nand2_x0 1 0 1675 1349 1352 nand2_x0
xsubckt_1008_nand3_x0 1 0 1328 1332 404 524 nand3_x0
xsubckt_507_a2_x2 0 171 1 233 538 a2_x2
xsubckt_459_a3_x2 1 218 0 219 220 221 a3_x2
xsubckt_449_a3_x2 1 228 0 229 234 235 a3_x2
xsubckt_224_nand4_x0 1 0 452 490 554 1730 591 nand4_x0
xsubckt_263_a2_x2 0 413 1 415 417 a2_x2
xsubckt_815_oa22_x2 0 1465 1 331 446 557 oa22_x2
xsubckt_1059_nand2_x0 1 0 1290 438 1724 nand2_x0
xsubckt_1227_oa22_x2 0 1146 1 1147 1173 656 oa22_x2
xsubckt_614_nand4_x0 1 0 69 551 552 554 1750 nand4_x0
xsubckt_1619_oa22_x2 0 787 1 24 956 789 oa22_x2
xsubckt_1396_nand3_x0 1 0 1006 383 554 1868 nand3_x0
xsubckt_1359_nand2_x0 1 0 1040 1130 1780 nand2_x0
xsubckt_580_nor4_x0 1 0 100 153 267 282 379 nor4_x0
xsubckt_221_nand2_x0 1 0 455 457 556 nand2_x0
xsubckt_723_oa22_x2 0 1549 1 281 360 626 oa22_x2
xsubckt_961_ao22_x2 0 1682 1 438 300 1367 ao22_x2
xsubckt_998_a3_x2 1 1338 0 516 520 538 a3_x2
xsubckt_1840_sff1_x4 1 9 0 1643 1766 sff1_x4
xsubckt_1801_sff1_x4 1 9 0 1674 1760 sff1_x4
xsubckt_1659_nand2_x0 1 0 747 749 925 nand2_x0
xsubckt_1332_a3_x2 1 1064 0 1065 1070 1078 a3_x2
xsubckt_485_nand3_x0 1 0 192 338 467 495 nand3_x0
xsubckt_235_oa22_x2 0 441 1 444 448 555 oa22_x2
xsubckt_700_o2_x2 0 1570 1 51 614 o2_x2
xsubckt_701_nand2_x0 1 0 1569 46 1848 nand2_x0
xsubckt_758_oa22_x2 0 1515 1 1521 1522 611 oa22_x2
xsubckt_1875_sff1_x4 1 9 0 1609 1779 sff1_x4
xsubckt_1527_oa22_x2 0 879 1 1561 956 881 oa22_x2
xsubckt_575_o2_x2 0 5 1 105 111 o2_x2
xsubckt_127_nand3_x0 1 0 549 551 552 554 nand3_x0
xsubckt_734_nand4_x0 1 0 1539 551 586 1725 1727 nand4_x0
xsubckt_918_ao22_x2 0 1379 1 1387 1383 1384 ao22_x2
xsubckt_1836_sff1_x4 1 9 0 1647 1790 sff1_x4
xsubckt_1440_a2_x2 0 965 1 966 968 a2_x2
xsubckt_1430_a2_x2 0 975 1 461 635 a2_x2
xsubckt_164_nand4_x0 1 0 512 516 521 527 532 nand4_x0
xsubckt_695_nand3_x0 1 0 1575 58 64 1840 nand3_x0
xsubckt_1135_mx2_x2 0 1643 1 1240 1232 1766 mx2_x2
xsubckt_1245_a2_x2 0 1144 1 546 550 a2_x2
xsubckt_1783_sff1_x4 1 9 0 1691 1825 sff1_x4
xsubckt_1579_a2_x2 0 827 1 828 831 a2_x2
xsubckt_1559_a2_x2 0 847 1 848 925 a2_x2
xsubckt_1483_mx2_x2 0 922 1 945 923 929 mx2_x2
xsubckt_1481_mx2_x2 0 924 1 930 927 940 mx2_x2
xsubckt_585_nor2_x0 1 0 96 305 396 nor2_x0
xsubckt_478_nand2_x0 1 0 199 200 539 nand2_x0
xsubckt_427_nand3_x0 1 0 250 415 417 420 nand3_x0
xsubckt_251_nand2_x0 1 0 425 481 495 nand2_x0
xsubckt_989_mx2_x2 0 1674 1 438 1348 1760 mx2_x2
xsubckt_1138_mx2_x2 0 1229 1 550 377 660 mx2_x2
xsubckt_958_nand2_x0 1 0 1683 1369 1371 nand2_x0
xsubckt_1779_sff1_x4 1 9 0 1695 1829 sff1_x4
xsubckt_1700_oa22_x2 0 706 1 709 711 739 oa22_x2
xsubckt_1372_nand2_x0 1 0 1028 1130 1779 nand2_x0
xsubckt_219_a4_x2 0 457 1 551 552 1726 587 a4_x2
xsubckt_778_nand2_x0 1 0 1497 1498 1503 nand2_x0
xsubckt_1621_nand3_x0 1 0 785 481 554 1774 nand3_x0
xsubckt_1368_nand3_x0 1 0 1031 1033 1042 1051 nand3_x0
xsubckt_444_a4_x2 0 233 1 528 530 534 536 a4_x2
xsubckt_93_inv_x0 1 0 1889 575 inv_x0
xsubckt_92_inv_x0 1 0 1810 576 inv_x0
xsubckt_91_inv_x0 1 0 1794 577 inv_x0
xsubckt_90_inv_x0 1 0 1890 578 inv_x0
xsubckt_229_a4_x2 0 447 1 1728 1727 1730 1729 a4_x2
xsubckt_1104_nand2_x0 1 0 1252 1253 1337 nand2_x0
xsubckt_1587_o2_x2 0 819 1 951 561 o2_x2
xsubckt_1411_ao22_x2 0 992 1 558 1138 993 ao22_x2
xsubckt_141_a2_x2 0 535 1 536 546 a2_x2
xsubckt_99_inv_x0 1 0 1887 569 inv_x0
xsubckt_98_inv_x0 1 0 1808 570 inv_x0
xsubckt_97_inv_x0 1 0 1792 571 inv_x0
xsubckt_96_inv_x0 1 0 1888 572 inv_x0
xsubckt_95_inv_x0 1 0 1809 573 inv_x0
xsubckt_94_inv_x0 1 0 1793 574 inv_x0
xsubckt_230_nand3_x0 1 0 446 447 586 1725 nand3_x0
xsubckt_289_a4_x2 0 387 1 476 587 1728 589 a4_x2
xsubckt_800_oa22_x2 0 1478 1 1521 1522 606 oa22_x2
xsubckt_851_nand2_x0 1 0 1902 1435 1439 nand2_x0
xsubckt_1137_nand4_x0 1 0 1230 473 495 585 641 nand4_x0
xsubckt_1170_nor2_x0 1 0 1201 1740 1759 nor2_x0
xsubckt_1682_oa22_x2 0 724 1 727 728 926 oa22_x2
xsubckt_1604_nxr2_x1 802 1 0 810 916 nxr2_x1
xsubckt_572_a3_x2 1 107 0 246 253 311 a3_x2
xsubckt_402_o4_x2 0 274 1 1728 1727 1730 1729 o4_x2
xsubckt_387_a3_x2 1 289 0 551 588 1727 a3_x2
xsubckt_154_ao22_x2 0 522 1 1786 1803 546 ao22_x2
xsubckt_151_a2_x2 0 525 1 527 532 a2_x2
xsubckt_161_a2_x2 0 515 1 516 521 a2_x2
xsubckt_171_a2_x2 0 505 1 508 510 a2_x2
xsubckt_181_a2_x2 0 495 1 586 1725 a2_x2
xsubckt_963_a4_x2 0 1365 1 404 439 525 539 a4_x2
xsubckt_640_a2_x2 0 43 1 44 343 a2_x2
xsubckt_530_nand3_x0 1 0 148 467 473 495 nand3_x0
xsubckt_403_nand2_x0 1 0 273 275 451 nand2_x0
xsubckt_856_a3_x2 1 1430 0 1431 1432 1433 a3_x2
xsubckt_1678_oa22_x2 0 728 1 734 736 939 oa22_x2
xsubckt_1354_ao22_x2 0 1044 1 563 1138 1045 ao22_x2
xsubckt_546_ao22_x2 0 133 1 327 188 134 ao22_x2
xsubckt_704_oa22_x2 0 1877 1 83 1571 1567 oa22_x2
xsubckt_769_a2_x2 0 1505 1 1506 1507 a2_x2
xsubckt_782_oa22_x2 0 1494 1 1521 1522 608 oa22_x2
xsubckt_1155_oa22_x2 0 1214 1 485 495 550 oa22_x2
xsubckt_1860_sff1_x4 1 9 0 1624 1869 sff1_x4
xsubckt_1821_sff1_x4 1 9 0 1654 1739 sff1_x4
xsubckt_133_nand2_x0 1 0 543 565 1786 nand2_x0
xsubckt_967_nand3_x0 1 0 1362 1365 150 413 nand3_x0
xsubckt_1005_a3_x2 1 1331 0 1360 412 538 a3_x2
xsubckt_1200_a3_x2 1 1173 0 1174 1181 1184 a3_x2
xsubckt_1720_mx2_x2 0 686 1 844 860 862 mx2_x2
xsubckt_1547_oa22_x2 0 859 1 911 864 906 oa22_x2
xsubckt_1514_a3_x2 1 892 0 932 937 1797 a3_x2
xsubckt_523_nand2_x0 1 0 155 457 467 nand2_x0
xsubckt_651_oa22_x2 0 33 1 281 360 632 oa22_x2
xsubckt_739_oa22_x2 0 1534 1 494 492 291 oa22_x2
xsubckt_1223_ao22_x2 0 1150 1 1173 1162 1151 ao22_x2
xsubckt_1262_ao22_x2 0 1127 1 1130 372 1782 ao22_x2
xsubckt_1856_sff1_x4 1 9 0 1628 1873 sff1_x4
xsubckt_1817_sff1_x4 1 9 0 1658 1732 sff1_x4
xsubckt_1723_mx2_x2 0 683 1 871 886 888 mx2_x2
xsubckt_1494_oa22_x2 0 911 1 1524 460 622 oa22_x2
xsubckt_1336_mx2_x2 0 1613 1 656 1061 1769 mx2_x2
xsubckt_1291_nand3_x0 1 0 1101 545 550 1862 nand3_x0
xsubckt_560_nand3_x0 1 0 119 289 467 493 nand3_x0
xsubckt_308_xr2_x1 368 0 1 1761 1855 xr2_x1
xsubckt_697_nand3_x0 1 0 1573 1574 1575 1576 nand3_x0
xsubckt_1644_nand2_x0 1 0 762 763 1046 nand2_x0
xsubckt_429_nand3_x0 1 0 248 251 504 538 nand3_x0
xsubckt_380_nand3_x0 1 0 296 467 481 554 nand3_x0
xsubckt_202_nand3_x0 1 0 474 476 490 554 nand3_x0
xsubckt_885_ao22_x2 0 1406 1 1409 1411 1852 ao22_x2
xsubckt_1258_ao22_x2 0 1131 1 1132 1135 1143 ao22_x2
xsubckt_1764_sff1_x4 1 9 0 1704 1814 sff1_x4
xsubckt_1298_mx2_x2 0 1617 1 656 1095 1773 mx2_x2
xsubckt_339_nand3_x0 1 0 337 490 590 1729 nand3_x0
xsubckt_1019_nand4_x0 1 0 1318 1322 1323 1344 1347 nand4_x0
xsubckt_1799_sff1_x4 1 9 0 1676 1735 sff1_x4
xsubckt_1523_ao22_x2 0 883 1 558 951 994 ao22_x2
xsubckt_1374_nand2_x0 1 0 1026 372 1850 nand2_x0
xsubckt_516_oa22_x2 0 162 1 163 185 555 oa22_x2
xsubckt_270_ao22_x2 0 406 1 511 507 420 ao22_x2
xsubckt_312_a4_x2 0 364 1 365 370 380 384 a4_x2
xsubckt_680_nand3_x0 1 0 1589 58 64 1841 nand3_x0
xsubckt_754_ao22_x2 0 1519 1 492 337 446 ao22_x2
xsubckt_1623_nand3_x0 1 0 783 932 937 1801 nand3_x0
xsubckt_1455_o2_x2 0 950 1 951 557 o2_x2
xsubckt_1284_nand2_x0 1 0 1107 1108 1113 nand2_x0
xsubckt_639_nand3_x0 1 0 44 338 495 1741 nand3_x0
xsubckt_616_a4_x2 0 67 1 273 320 334 336 a4_x2
xsubckt_372_a4_x2 0 304 1 306 329 340 363 a4_x2
xsubckt_196_nand4_x0 1 0 480 1728 589 1730 591 nand4_x0
xsubckt_1716_oa22_x2 0 690 1 841 826 823 oa22_x2
xsubckt_1470_ao22_x2 0 935 1 494 480 309 ao22_x2
xsubckt_420_a3_x2 1 257 0 413 504 538 a3_x2
xsubckt_283_nand2_x0 1 0 393 394 395 nand2_x0
xsubckt_820_oa22_x2 0 1893 1 1550 1543 1461 oa22_x2
xsubckt_853_nand2_x0 1 0 1433 1458 1868 nand2_x0
xsubckt_871_a4_x2 0 1419 1 551 552 554 660 a4_x2
xsubckt_908_oa22_x2 0 1387 1 1389 1391 645 oa22_x2
xsubckt_980_nand3_x0 1 0 1353 1365 406 413 nand3_x0
xsubckt_1406_nand2_x0 1 0 997 1130 1776 nand2_x0
xsubckt_490_a3_x2 1 187 0 189 198 201 a3_x2
xsubckt_371_oa22_x2 0 305 1 1723 442 308 oa22_x2
xsubckt_135_ao22_x2 0 541 1 1786 1799 546 ao22_x2
xsubckt_228_nand4_x0 1 0 448 451 490 1730 591 nand4_x0
xsubckt_303_a2_x2 0 373 1 374 376 a2_x2
xsubckt_313_a2_x2 0 363 1 364 373 a2_x2
xsubckt_1049_nand4_x0 1 0 1297 1332 404 439 525 nand4_x0
xsubckt_1427_ao22_x2 0 978 1 1523 461 1733 ao22_x2
xsubckt_617_a2_x2 0 66 1 67 69 a2_x2
xsubckt_589_a3_x2 1 92 0 210 347 462 a3_x2
xsubckt_383_a2_x2 0 293 1 294 296 a2_x2
xsubckt_373_a2_x2 0 303 1 304 311 a2_x2
xsubckt_168_a2_x2 0 508 1 509 546 a2_x2
xsubckt_669_nand3_x0 1 0 17 58 64 1842 nand3_x0
xsubckt_794_a3_x2 1 1483 0 1484 1487 1488 a3_x2
xsubckt_816_oa22_x2 0 1464 1 1521 1522 604 oa22_x2
xsubckt_1140_oa22_x2 0 1227 1 239 1229 1231 oa22_x2
xsubckt_527_ao22_x2 0 151 1 243 236 152 ao22_x2
xsubckt_442_nand3_x0 1 0 235 244 432 478 nand3_x0
xsubckt_352_nand3_x0 1 0 324 447 467 554 nand3_x0
xsubckt_724_oa22_x2 0 1548 1 44 343 636 oa22_x2
xsubckt_763_oa22_x2 0 1906 1 52 1543 1511 oa22_x2
xsubckt_973_nand2_x0 1 0 1358 438 1736 nand2_x0
xsubckt_1880_sff1_x4 1 9 0 1604 1856 sff1_x4
xsubckt_1731_ao22_x2 0 675 1 676 677 700 ao22_x2
xsubckt_1364_a4_x2 0 1035 1 1036 1037 1038 343 a4_x2
xsubckt_489_nand3_x0 1 0 188 437 541 543 nand3_x0
xsubckt_348_nand4_x0 1 0 328 447 467 586 1725 nand4_x0
xsubckt_341_o2_x2 0 335 1 336 555 o2_x2
xsubckt_166_o2_x2 0 510 1 1796 1786 o2_x2
xsubckt_1841_sff1_x4 1 9 0 1642 1795 sff1_x4
xsubckt_1802_sff1_x4 1 9 0 1673 1745 sff1_x4
xsubckt_525_nand2_x0 1 0 153 155 156 nand2_x0
xsubckt_511_nand4_x0 1 0 167 517 520 527 532 nand4_x0
xsubckt_236_oa22_x2 0 440 1 662 442 459 oa22_x2
xsubckt_759_oa22_x2 0 1514 1 331 446 564 oa22_x2
xsubckt_1876_sff1_x4 1 9 0 1608 1778 sff1_x4
xsubckt_1837_sff1_x4 1 9 0 1646 1789 sff1_x4
xsubckt_1520_a2_x2 0 886 1 887 905 a2_x2
xsubckt_1510_a2_x2 0 896 1 897 978 a2_x2
xsubckt_1335_a2_x2 0 1061 1 1062 1063 a2_x2
xsubckt_255_mx2_x2 0 421 1 1786 1797 1788 mx2_x2
xsubckt_675_o2_x2 0 11 1 51 617 o2_x2
xsubckt_789_nand3_x0 1 0 1488 1518 1526 1772 nand3_x0
xsubckt_1071_a2_x2 0 1280 1 1281 1330 a2_x2
xsubckt_1081_a2_x2 0 1271 1 1329 439 a2_x2
xsubckt_1629_a2_x2 0 777 1 778 925 a2_x2
xsubckt_1436_oa22_x2 0 969 1 970 972 1738 oa22_x2
xsubckt_1365_a2_x2 0 1034 1 1035 1039 a2_x2
xsubckt_1355_a2_x2 0 1043 1 1044 1049 a2_x2
xsubckt_345_nand2_x0 1 0 331 338 493 nand2_x0
xsubckt_331_nand4_x0 1 0 345 476 554 588 1727 nand4_x0
xsubckt_204_nand3_x0 1 0 472 551 1728 589 nand3_x0
xsubckt_667_oa22_x2 0 1880 1 83 24 19 oa22_x2
xsubckt_1146_mx2_x2 0 1222 1 549 1223 377 mx2_x2
xsubckt_1147_mx2_x2 0 1221 1 660 1850 653 mx2_x2
xsubckt_1148_mx2_x2 0 1220 1 378 1221 1800 mx2_x2
xsubckt_1149_mx2_x2 0 1641 1 1222 1220 1812 mx2_x2
xsubckt_1784_sff1_x4 1 9 0 1690 1824 sff1_x4
xsubckt_1740_nxr2_x1 671 1 0 689 692 nxr2_x1
xsubckt_1689_a2_x2 0 717 1 718 963 a2_x2
xsubckt_1466_nand2_x0 1 0 939 941 943 nand2_x0
xsubckt_378_nand4_x0 1 0 298 404 409 437 525 nand4_x0
xsubckt_292_nand3_x0 1 0 384 387 467 1726 nand3_x0
xsubckt_772_nand3_x0 1 0 1503 1518 1526 1774 nand3_x0
xsubckt_1582_ao22_x2 0 824 1 835 837 915 ao22_x2
xsubckt_1490_o3_x2 0 915 1 918 919 84 o3_x2
xsubckt_1305_oa22_x2 0 1088 1 1772 1128 1090 oa22_x2
xsubckt_631_nand4_x0 1 0 52 53 54 55 56 nand4_x0
xsubckt_682_nand3_x0 1 0 1587 58 63 1825 nand3_x0
xsubckt_1162_nor4_x0 1 0 1208 1846 1847 1848 1849 nor4_x0
xsubckt_1617_o2_x2 0 789 1 791 793 o2_x2
xsubckt_678_nand4_x0 1 0 1590 1591 10 11 12 nand4_x0
xsubckt_1108_nand2_x0 1 0 1248 1249 1251 nand2_x0
xsubckt_1578_ao22_x2 0 828 1 829 838 977 ao22_x2
xsubckt_612_a3_x2 1 71 0 72 75 241 a3_x2
xsubckt_407_a3_x2 1 269 0 275 1726 587 a3_x2
xsubckt_361_nand4_x0 1 0 315 447 467 1726 587 nand4_x0
xsubckt_173_a3_x2 1 503 0 505 520 532 a3_x2
xsubckt_208_ao22_x2 0 468 1 472 492 1723 ao22_x2
xsubckt_855_nand2_x0 1 0 1431 1531 1798 nand2_x0
xsubckt_1018_nand2_x0 1 0 1319 438 624 nand2_x0
xsubckt_1145_nor3_x0 1 0 1223 1736 1758 1740 nor3_x0
xsubckt_1616_nor2_x0 1 0 790 791 793 nor2_x0
xsubckt_1486_ao22_x2 0 919 1 1523 461 1743 ao22_x2
xsubckt_1408_nand2_x0 1 0 995 372 1847 nand2_x0
xsubckt_1287_oa22_x2 0 1104 1 1124 1115 1107 oa22_x2
xsubckt_624_nand3_x0 1 0 59 61 71 77 nand3_x0
xsubckt_505_a2_x2 0 173 1 517 520 a2_x2
xsubckt_487_a3_x2 1 190 0 191 192 193 a3_x2
xsubckt_261_a2_x2 0 415 1 416 546 a2_x2
xsubckt_565_a2_x2 0 114 1 115 116 a2_x2
xsubckt_535_a2_x2 0 143 1 144 146 a2_x2
xsubckt_497_a3_x2 1 181 0 182 184 254 a3_x2
xsubckt_309_nxr2_x1 367 1 0 1761 1855 nxr2_x1
xsubckt_661_nand4_x0 1 0 24 26 27 28 29 nand4_x0
xsubckt_692_a3_x2 1 1578 0 58 63 1824 a3_x2
xsubckt_1001_nand2_x0 1 0 1335 412 505 nand2_x0
xsubckt_1160_oa22_x2 0 1210 1 389 495 1740 oa22_x2
xsubckt_1591_oa22_x2 0 815 1 1850 952 817 oa22_x2
xsubckt_783_oa22_x2 0 1493 1 331 446 561 oa22_x2
xsubckt_975_nand2_x0 1 0 1678 1357 1358 nand2_x0
xsubckt_1552_oa22_x2 0 854 1 1848 952 856 oa22_x2
xsubckt_1301_nand2_x0 1 0 1092 1094 343 nand2_x0
xsubckt_104_mx2_x2 0 564 1 656 578 579 mx2_x2
xsubckt_834_nand3_x0 1 0 1449 1518 1526 1780 nand3_x0
xsubckt_1861_sff1_x4 1 9 0 1623 1868 sff1_x4
xsubckt_1822_sff1_x4 1 9 0 1803 1811 sff1_x4
xsubckt_108_mx2_x2 0 562 1 656 572 573 mx2_x2
xsubckt_106_mx2_x2 0 563 1 656 575 576 mx2_x2
xsubckt_652_oa22_x2 0 32 1 48 482 651 oa22_x2
xsubckt_691_oa22_x2 0 1878 1 83 1584 1579 oa22_x2
xsubckt_779_oa22_x2 0 1898 1 24 1543 1497 oa22_x2
xsubckt_795_nand2_x0 1 0 1896 1483 1489 nand2_x0
xsubckt_1857_sff1_x4 1 9 0 1627 1872 sff1_x4
xsubckt_1818_sff1_x4 1 9 0 1657 1731 sff1_x4
xsubckt_1509_oa22_x2 0 897 1 52 956 898 oa22_x2
xsubckt_1479_a3_x2 1 926 0 928 941 943 a3_x2
xsubckt_1385_nand3_x0 1 0 1016 383 554 1869 nand3_x0
xsubckt_564_nand3_x0 1 0 115 389 495 556 nand3_x0
xsubckt_398_o2_x2 0 278 1 279 555 o2_x2
xsubckt_1099_oa22_x2 0 1654 1 1739 549 2 oa22_x2
xsubckt_1213_a2_x2 0 1160 1 386 446 a2_x2
xsubckt_1739_mx2_x2 0 1599 1 656 702 1850 mx2_x2
xsubckt_1738_mx2_x2 0 1600 1 656 696 1851 mx2_x2
xsubckt_1737_mx2_x2 0 1601 1 656 698 1852 mx2_x2
xsubckt_1736_mx2_x2 0 1602 1 656 672 1853 mx2_x2
xsubckt_1722_a2_x2 0 684 1 871 887 a2_x2
xsubckt_1694_ao22_x2 0 712 1 715 716 720 ao22_x2
xsubckt_1348_mx2_x2 0 1612 1 656 1050 1768 mx2_x2
xsubckt_600_nand2_x0 1 0 82 489 494 nand2_x0
xsubckt_474_nand3_x0 1 0 203 402 515 539 nand3_x0
xsubckt_827_nand2_x0 1 0 1892 1455 1460 nand2_x0
xsubckt_1078_nand2_x0 1 0 1274 438 581 nand2_x0
xsubckt_1765_sff1_x4 1 9 0 8 1730 sff1_x4
xsubckt_1655_ao22_x2 0 751 1 755 757 940 ao22_x2
xsubckt_1595_nand3_x0 1 0 811 932 937 1800 nand3_x0
xsubckt_1577_a2_x2 0 829 1 830 925 a2_x2
xsubckt_1558_nand2_x0 1 0 848 849 850 nand2_x0
xsubckt_510_nand2_x0 1 0 168 232 249 nand2_x0
xsubckt_167_nand2_x0 1 0 509 598 1786 nand2_x0
xsubckt_257_nand2_x0 1 0 419 421 546 nand2_x0
xsubckt_864_nand3_x0 1 0 1424 1518 1526 1775 nand3_x0
xsubckt_1698_mx2_x2 0 708 1 743 740 741 mx2_x2
xsubckt_1325_oa22_x2 0 1070 1 1770 1128 1072 oa22_x2
xsubckt_227_a4_x2 0 449 1 451 490 1730 591 a4_x2
xsubckt_237_a4_x2 0 439 1 551 552 554 1721 a4_x2
xsubckt_240_nand2_x0 1 0 436 439 655 nand2_x0
xsubckt_909_nxr2_x1 1386 1 0 1388 1848 nxr2_x1
xsubckt_326_nand3_x0 1 0 350 362 467 495 nand3_x0
xsubckt_150_nand2_x0 1 0 526 529 531 nand2_x0
xsubckt_806_nand3_x0 1 0 1473 1518 1526 1770 nand3_x0
xsubckt_857_nand2_x0 1 0 1901 1430 1434 nand2_x0
xsubckt_984_nand3_x0 1 0 1350 419 506 509 nand3_x0
xsubckt_1094_nand4_x0 1 0 1260 1351 413 517 520 nand4_x0
xsubckt_1664_nxr2_x1 742 1 0 753 915 nxr2_x1
xsubckt_540_a3_x2 1 138 0 139 318 326 a3_x2
xsubckt_365_a3_x2 1 311 0 312 318 326 a3_x2
xsubckt_197_nand2_x0 1 0 479 481 493 nand2_x0
xsubckt_991_a4_x2 0 1345 1 420 504 517 520 a4_x2
xsubckt_1220_nand3_x0 1 0 1153 1169 1534 82 nand3_x0
xsubckt_453_a2_x2 0 224 1 225 227 a2_x2
xsubckt_844_a3_x2 1 1440 0 1441 1442 1443 a3_x2
xsubckt_1130_nand3_x0 1 0 1236 1237 1419 654 nand3_x0
xsubckt_1141_oa22_x2 0 1226 1 1228 1230 668 oa22_x2
xsubckt_1180_oa22_x2 0 1193 1 288 472 492 oa22_x2
xsubckt_446_nand3_x0 1 0 231 233 516 520 nand3_x0
xsubckt_280_oa22_x2 0 396 1 437 399 424 oa22_x2
xsubckt_285_o4_x2 0 391 1 393 428 433 440 o4_x2
xsubckt_298_a2_x2 0 378 1 389 495 a2_x2
xsubckt_305_nand4_x0 1 0 371 476 554 1728 589 nand4_x0
xsubckt_1091_nand2_x0 1 0 1262 1263 1368 nand2_x0
xsubckt_1533_oa22_x2 0 873 1 876 877 926 oa22_x2
xsubckt_1414_a4_x2 0 989 1 990 1002 1011 1020 a4_x2
xsubckt_1340_nand3_x0 1 0 1057 383 554 1873 nand3_x0
xsubckt_528_ao22_x2 0 150 1 511 507 419 ao22_x2
xsubckt_209_nor2_x0 1 0 467 2 1721 nor2_x0
xsubckt_725_oa22_x2 0 1547 1 48 482 642 oa22_x2
xsubckt_746_nand3_x0 1 0 1527 1528 1530 1532 nand3_x0
xsubckt_1881_sff1_x4 1 9 0 1603 1855 sff1_x4
xsubckt_1842_sff1_x4 1 9 0 1641 1812 sff1_x4
xsubckt_1803_sff1_x4 1 9 0 1672 1744 sff1_x4
xsubckt_1512_a3_x2 1 894 0 481 554 1770 a3_x2
xsubckt_656_nand3_x0 1 0 29 57 63 1819 nand3_x0
xsubckt_799_oa22_x2 0 1479 1 331 446 559 oa22_x2
xsubckt_1111_a2_x2 0 1246 1 193 313 a2_x2
xsubckt_1123_nand2_x0 1 0 1243 461 1760 nand2_x0
xsubckt_1877_sff1_x4 1 9 0 1607 1777 sff1_x4
xsubckt_1610_a2_x2 0 796 1 800 804 a2_x2
xsubckt_1600_a2_x2 0 806 1 807 925 a2_x2
xsubckt_1529_oa22_x2 0 877 1 891 893 939 oa22_x2
xsubckt_1367_a3_x2 1 1032 0 1033 1042 1051 a3_x2
xsubckt_1283_ao22_x2 0 1108 1 648 1136 1109 ao22_x2
xsubckt_515_nand4_x0 1 0 163 164 169 178 181 nand4_x0
xsubckt_1205_ao22_x2 0 1168 1 292 481 554 ao22_x2
xsubckt_1838_sff1_x4 1 9 0 1645 1788 sff1_x4
xsubckt_1750_sff1_x4 1 9 0 1718 1844 sff1_x4
xsubckt_1719_a2_x2 0 687 1 844 861 a2_x2
xsubckt_1476_oa22_x2 0 929 1 931 938 939 oa22_x2
xsubckt_1465_a2_x2 0 940 1 941 943 a2_x2
xsubckt_602_nand2_x0 1 0 80 81 1724 nand2_x0
xsubckt_386_nand3_x0 1 0 290 292 467 495 nand3_x0
xsubckt_349_nand2_x0 1 0 327 526 533 nand2_x0
xsubckt_829_nand2_x0 1 0 1453 1458 1872 nand2_x0
xsubckt_1011_o3_x2 0 1325 1 1327 1333 1339 o3_x2
xsubckt_1070_nand3_x0 1 0 1281 1351 412 533 nand3_x0
xsubckt_1156_mx2_x2 0 1213 1 1214 1796 1846 mx2_x2
xsubckt_1785_sff1_x4 1 9 0 1689 1823 sff1_x4
xsubckt_1437_oa22_x2 0 968 1 369 471 644 oa22_x2
xsubckt_169_nand2_x0 1 0 507 509 546 nand2_x0
xsubckt_296_nand3_x0 1 0 380 383 493 556 nand3_x0
xsubckt_740_ao22_x2 0 1533 1 495 493 292 ao22_x2
xsubckt_1152_ao22_x2 0 1217 1 58 63 1746 ao22_x2
xsubckt_1157_mx2_x2 0 1640 1 1215 1785 1213 mx2_x2
xsubckt_1153_nand2_x0 1 0 1216 1419 657 nand2_x0
xsubckt_1228_o2_x2 0 1145 1 1146 1150 o2_x2
xsubckt_1670_nand3_x0 1 0 736 481 554 1782 nand3_x0
xsubckt_1505_ao22_x2 0 901 1 954 1540 1853 ao22_x2
xsubckt_455_nand4_x0 1 0 222 402 437 515 538 nand4_x0
xsubckt_332_nand2_x0 1 0 344 346 467 nand2_x0
xsubckt_330_a4_x2 0 346 1 476 554 588 1727 a4_x2
xsubckt_203_a3_x2 1 473 0 551 1728 589 a3_x2
xsubckt_812_nand2_x0 1 0 1894 1468 1474 nand2_x0
xsubckt_990_nand2_x0 1 0 1346 438 625 nand2_x0
xsubckt_1163_nor4_x0 1 0 1207 1850 1851 1852 1853 nor4_x0
xsubckt_1453_nand2_x0 1 0 952 955 1541 nand2_x0
xsubckt_1402_nand3_x0 1 0 1000 1002 1011 1020 nand3_x0
xsubckt_379_nand2_x0 1 0 297 481 554 nand2_x0
xsubckt_328_nand3_x0 1 0 348 358 495 556 nand3_x0
xsubckt_152_nand2_x0 1 0 524 527 532 nand2_x0
xsubckt_195_a4_x2 0 481 1 1728 589 1730 591 a4_x2
xsubckt_859_nand2_x0 1 0 1428 1458 1867 nand2_x0
xsubckt_1363_nand2_x0 1 0 1036 372 1851 nand2_x0
xsubckt_628_nand3_x0 1 0 55 57 63 1821 nand3_x0
xsubckt_557_a3_x2 1 122 0 123 130 133 a3_x2
xsubckt_321_a2_x2 0 355 1 358 493 a2_x2
xsubckt_684_a4_x2 0 1585 1 1586 1587 1588 1589 a4_x2
xsubckt_718_nand3_x0 1 0 1554 57 64 1830 nand3_x0
xsubckt_732_a3_x2 1 1541 0 1542 351 375 a3_x2
xsubckt_1017_ao22_x2 0 1673 1 1321 1324 1346 ao22_x2
xsubckt_615_a2_x2 0 68 1 273 336 a2_x2
xsubckt_538_nand3_x0 1 0 140 467 473 493 nand3_x0
xsubckt_362_nand2_x0 1 0 314 323 1726 nand2_x0
xsubckt_311_nand3_x0 1 0 365 366 383 554 nand3_x0
xsubckt_752_a3_x2 1 1521 0 371 445 479 a3_x2
xsubckt_810_a2_x2 0 1469 1 1470 1471 a2_x2
xsubckt_1183_nand2_x0 1 0 1190 1193 1194 nand2_x0
xsubckt_1573_nand2_x0 1 0 833 834 836 nand2_x0
xsubckt_499_nand2_x0 1 0 179 180 400 nand2_x0
xsubckt_448_nand3_x0 1 0 229 232 405 437 nand3_x0
xsubckt_842_nand2_x0 1 0 1442 1531 1800 nand2_x0
xsubckt_870_a2_x2 0 1592 1 1763 1812 a2_x2
xsubckt_979_nand2_x0 1 0 1354 438 1735 nand2_x0
xsubckt_1179_nand3_x0 1 0 1194 551 554 1728 nand3_x0
xsubckt_1342_a4_x2 0 1055 1 1056 1057 1058 343 a4_x2
xsubckt_509_ao22_x2 0 169 1 231 176 170 ao22_x2
xsubckt_110_mx2_x2 0 561 1 656 569 570 mx2_x2
xsubckt_182_nand2_x0 1 0 494 586 1725 nand2_x0
xsubckt_268_nand3_x0 1 0 408 412 504 538 nand3_x0
xsubckt_959_a2_x2 0 1368 1 299 439 a2_x2
xsubckt_1862_sff1_x4 1 9 0 1622 1867 sff1_x4
xsubckt_1823_sff1_x4 1 9 0 1802 1810 sff1_x4
xsubckt_1713_ao22_x2 0 693 1 703 796 797 ao22_x2
xsubckt_1393_nand2_x0 1 0 1009 1130 1777 nand2_x0
xsubckt_633_o2_x2 0 50 1 51 620 o2_x2
xsubckt_116_mx2_x2 0 558 1 656 596 597 mx2_x2
xsubckt_114_mx2_x2 0 559 1 656 593 594 mx2_x2
xsubckt_112_mx2_x2 0 560 1 656 566 567 mx2_x2
xsubckt_178_nand3_x0 1 0 498 552 1730 591 nand3_x0
xsubckt_658_nand3_x0 1 0 27 57 64 1835 nand3_x0
xsubckt_1252_nand3_x0 1 0 1137 1534 385 491 nand3_x0
.ends Arlet6502
